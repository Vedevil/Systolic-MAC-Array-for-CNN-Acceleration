magic
tech sky130A
magscale 1 2
timestamp 1760531949
<< viali >>
rect 7389 16609 7423 16643
rect 7481 16609 7515 16643
rect 7849 16609 7883 16643
rect 8401 16609 8435 16643
rect 11897 16609 11931 16643
rect 12081 16609 12115 16643
rect 5365 16541 5399 16575
rect 7573 16541 7607 16575
rect 7665 16541 7699 16575
rect 11805 16541 11839 16575
rect 11989 16541 12023 16575
rect 4813 16405 4847 16439
rect 7205 16405 7239 16439
rect 11621 16405 11655 16439
rect 4997 16201 5031 16235
rect 9689 16201 9723 16235
rect 11253 16133 11287 16167
rect 12357 16133 12391 16167
rect 7113 16065 7147 16099
rect 10885 16065 10919 16099
rect 11345 16065 11379 16099
rect 12909 16065 12943 16099
rect 3249 15997 3283 16031
rect 3525 15997 3559 16031
rect 5641 15997 5675 16031
rect 7941 15997 7975 16031
rect 8217 15997 8251 16031
rect 11069 15997 11103 16031
rect 11529 15997 11563 16031
rect 5089 15861 5123 15895
rect 7665 15861 7699 15895
rect 12173 15861 12207 15895
rect 4892 15657 4926 15691
rect 7953 15657 7987 15691
rect 8309 15657 8343 15691
rect 13277 15657 13311 15691
rect 1869 15521 1903 15555
rect 4629 15521 4663 15555
rect 8217 15521 8251 15555
rect 10149 15521 10183 15555
rect 11805 15521 11839 15555
rect 3801 15453 3835 15487
rect 8493 15453 8527 15487
rect 9873 15453 9907 15487
rect 9965 15453 9999 15487
rect 10241 15453 10275 15487
rect 10701 15453 10735 15487
rect 11345 15453 11379 15487
rect 11529 15453 11563 15487
rect 13553 15453 13587 15487
rect 2145 15385 2179 15419
rect 3617 15317 3651 15351
rect 4445 15317 4479 15351
rect 6377 15317 6411 15351
rect 6469 15317 6503 15351
rect 9689 15317 9723 15351
rect 13461 15317 13495 15351
rect 3893 15113 3927 15147
rect 6929 15113 6963 15147
rect 7205 15113 7239 15147
rect 8309 15113 8343 15147
rect 8769 15113 8803 15147
rect 9229 15113 9263 15147
rect 7046 15045 7080 15079
rect 9689 15045 9723 15079
rect 2973 14977 3007 15011
rect 3249 14977 3283 15011
rect 3433 14977 3467 15011
rect 4077 14977 4111 15011
rect 4261 14977 4295 15011
rect 4445 14977 4479 15011
rect 6561 14977 6595 15011
rect 8401 14977 8435 15011
rect 9137 14977 9171 15011
rect 2697 14909 2731 14943
rect 3341 14909 3375 14943
rect 4353 14909 4387 14943
rect 4721 14909 4755 14943
rect 6837 14909 6871 14943
rect 7849 14909 7883 14943
rect 8217 14909 8251 14943
rect 9413 14909 9447 14943
rect 11989 14909 12023 14943
rect 12265 14909 12299 14943
rect 15301 14909 15335 14943
rect 15577 14909 15611 14943
rect 2789 14841 2823 14875
rect 2881 14773 2915 14807
rect 6193 14773 6227 14807
rect 7297 14773 7331 14807
rect 11161 14773 11195 14807
rect 13737 14773 13771 14807
rect 13829 14773 13863 14807
rect 4813 14569 4847 14603
rect 5457 14569 5491 14603
rect 8309 14569 8343 14603
rect 11713 14569 11747 14603
rect 12265 14569 12299 14603
rect 14749 14569 14783 14603
rect 5089 14501 5123 14535
rect 5641 14501 5675 14535
rect 13737 14501 13771 14535
rect 6285 14433 6319 14467
rect 6469 14433 6503 14467
rect 7021 14433 7055 14467
rect 7757 14433 7791 14467
rect 9137 14433 9171 14467
rect 12173 14433 12207 14467
rect 14565 14433 14599 14467
rect 4997 14365 5031 14399
rect 5273 14365 5307 14399
rect 5549 14365 5583 14399
rect 7297 14365 7331 14399
rect 7849 14365 7883 14399
rect 8125 14365 8159 14399
rect 8217 14365 8251 14399
rect 8401 14365 8435 14399
rect 10977 14365 11011 14399
rect 11161 14365 11195 14399
rect 11621 14365 11655 14399
rect 11989 14365 12023 14399
rect 12449 14365 12483 14399
rect 12541 14365 12575 14399
rect 13093 14365 13127 14399
rect 13277 14365 13311 14399
rect 13369 14365 13403 14399
rect 13553 14365 13587 14399
rect 13645 14365 13679 14399
rect 14473 14365 14507 14399
rect 15393 14365 15427 14399
rect 8033 14297 8067 14331
rect 9413 14297 9447 14331
rect 13461 14297 13495 14331
rect 14105 14297 14139 14331
rect 6009 14229 6043 14263
rect 6101 14229 6135 14263
rect 7297 14229 7331 14263
rect 7941 14229 7975 14263
rect 10885 14229 10919 14263
rect 11069 14229 11103 14263
rect 12909 14229 12943 14263
rect 13093 14229 13127 14263
rect 14841 14229 14875 14263
rect 5365 14025 5399 14059
rect 5457 14025 5491 14059
rect 9689 14025 9723 14059
rect 11161 14025 11195 14059
rect 2697 13889 2731 13923
rect 5089 13889 5123 13923
rect 5549 13889 5583 13923
rect 9413 13889 9447 13923
rect 9597 13889 9631 13923
rect 10609 13889 10643 13923
rect 13737 13889 13771 13923
rect 2881 13821 2915 13855
rect 2973 13821 3007 13855
rect 3341 13821 3375 13855
rect 3893 13821 3927 13855
rect 9045 13821 9079 13855
rect 9137 13821 9171 13855
rect 10333 13821 10367 13855
rect 13093 13821 13127 13855
rect 13645 13821 13679 13855
rect 14013 13821 14047 13855
rect 15485 13821 15519 13855
rect 2513 13685 2547 13719
rect 11069 13481 11103 13515
rect 13369 13481 13403 13515
rect 2053 13345 2087 13379
rect 8769 13345 8803 13379
rect 10333 13345 10367 13379
rect 10793 13345 10827 13379
rect 10885 13345 10919 13379
rect 13185 13345 13219 13379
rect 14105 13345 14139 13379
rect 14473 13345 14507 13379
rect 14565 13345 14599 13379
rect 1777 13277 1811 13311
rect 3801 13277 3835 13311
rect 4353 13277 4387 13311
rect 7021 13277 7055 13311
rect 9781 13277 9815 13311
rect 10425 13277 10459 13311
rect 10517 13277 10551 13311
rect 10609 13277 10643 13311
rect 11345 13277 11379 13311
rect 13645 13277 13679 13311
rect 14289 13277 14323 13311
rect 14381 13277 14415 13311
rect 7297 13209 7331 13243
rect 11253 13209 11287 13243
rect 13553 13209 13587 13243
rect 3525 13141 3559 13175
rect 9229 13141 9263 13175
rect 3617 12937 3651 12971
rect 5181 12937 5215 12971
rect 7757 12937 7791 12971
rect 5273 12869 5307 12903
rect 8309 12869 8343 12903
rect 9137 12869 9171 12903
rect 13645 12869 13679 12903
rect 4353 12801 4387 12835
rect 4629 12801 4663 12835
rect 4813 12801 4847 12835
rect 5181 12801 5215 12835
rect 5457 12801 5491 12835
rect 5733 12801 5767 12835
rect 6009 12801 6043 12835
rect 6193 12801 6227 12835
rect 7941 12801 7975 12835
rect 8585 12801 8619 12835
rect 10977 12801 11011 12835
rect 11069 12801 11103 12835
rect 13277 12801 13311 12835
rect 13737 12801 13771 12835
rect 13921 12801 13955 12835
rect 1869 12733 1903 12767
rect 2145 12733 2179 12767
rect 4169 12733 4203 12767
rect 8125 12733 8159 12767
rect 8217 12733 8251 12767
rect 8309 12733 8343 12767
rect 8861 12733 8895 12767
rect 10885 12733 10919 12767
rect 11161 12733 11195 12767
rect 12817 12733 12851 12767
rect 13185 12733 13219 12767
rect 5549 12597 5583 12631
rect 8493 12597 8527 12631
rect 10609 12597 10643 12631
rect 10701 12597 10735 12631
rect 12173 12597 12207 12631
rect 13553 12597 13587 12631
rect 13829 12597 13863 12631
rect 6561 12393 6595 12427
rect 9781 12393 9815 12427
rect 9965 12393 9999 12427
rect 13645 12393 13679 12427
rect 6653 12325 6687 12359
rect 9229 12325 9263 12359
rect 13093 12325 13127 12359
rect 3617 12257 3651 12291
rect 3985 12257 4019 12291
rect 8033 12257 8067 12291
rect 9873 12257 9907 12291
rect 10517 12257 10551 12291
rect 10793 12257 10827 12291
rect 1869 12189 1903 12223
rect 5273 12189 5307 12223
rect 6193 12189 6227 12223
rect 6561 12189 6595 12223
rect 7573 12189 7607 12223
rect 7665 12189 7699 12223
rect 8309 12189 8343 12223
rect 8493 12189 8527 12223
rect 9354 12189 9388 12223
rect 11161 12189 11195 12223
rect 11253 12189 11287 12223
rect 11345 12189 11379 12223
rect 13369 12189 13403 12223
rect 13461 12189 13495 12223
rect 13737 12189 13771 12223
rect 14197 12189 14231 12223
rect 14749 12189 14783 12223
rect 2145 12121 2179 12155
rect 6837 12121 6871 12155
rect 7757 12121 7791 12155
rect 7941 12121 7975 12155
rect 11621 12121 11655 12155
rect 4629 12053 4663 12087
rect 4721 12053 4755 12087
rect 5549 12053 5583 12087
rect 6929 12053 6963 12087
rect 9413 12053 9447 12087
rect 11069 12053 11103 12087
rect 13185 12053 13219 12087
rect 2421 11849 2455 11883
rect 6193 11849 6227 11883
rect 8217 11849 8251 11883
rect 10057 11849 10091 11883
rect 8309 11781 8343 11815
rect 13093 11781 13127 11815
rect 2605 11713 2639 11747
rect 2881 11713 2915 11747
rect 3801 11713 3835 11747
rect 4445 11713 4479 11747
rect 8493 11713 8527 11747
rect 8677 11713 8711 11747
rect 10149 11713 10183 11747
rect 11897 11713 11931 11747
rect 12817 11713 12851 11747
rect 3249 11645 3283 11679
rect 4077 11645 4111 11679
rect 4721 11645 4755 11679
rect 6469 11645 6503 11679
rect 6745 11645 6779 11679
rect 11529 11645 11563 11679
rect 12081 11645 12115 11679
rect 14565 11645 14599 11679
rect 3525 11577 3559 11611
rect 3709 11577 3743 11611
rect 8585 11577 8619 11611
rect 11621 11577 11655 11611
rect 2789 11509 2823 11543
rect 4169 11509 4203 11543
rect 4353 11509 4387 11543
rect 3893 11305 3927 11339
rect 4261 11305 4295 11339
rect 4537 11305 4571 11339
rect 4905 11305 4939 11339
rect 5444 11305 5478 11339
rect 7757 11305 7791 11339
rect 8033 11237 8067 11271
rect 13829 11237 13863 11271
rect 2973 11169 3007 11203
rect 3525 11169 3559 11203
rect 3617 11169 3651 11203
rect 4077 11169 4111 11203
rect 4445 11169 4479 11203
rect 4813 11169 4847 11203
rect 5181 11169 5215 11203
rect 8125 11169 8159 11203
rect 8217 11169 8251 11203
rect 9689 11169 9723 11203
rect 9965 11169 9999 11203
rect 11437 11169 11471 11203
rect 11805 11169 11839 11203
rect 12541 11169 12575 11203
rect 14473 11169 14507 11203
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 3341 11101 3375 11135
rect 3801 11101 3835 11135
rect 4353 11101 4387 11135
rect 4629 11101 4663 11135
rect 4721 11101 4755 11135
rect 4997 11101 5031 11135
rect 5089 11101 5123 11135
rect 7941 11101 7975 11135
rect 8401 11101 8435 11135
rect 8953 11101 8987 11135
rect 9505 11101 9539 11135
rect 12725 11101 12759 11135
rect 12817 11101 12851 11135
rect 13461 11101 13495 11135
rect 13645 11101 13679 11135
rect 13897 11101 13931 11135
rect 14565 11101 14599 11135
rect 3157 11033 3191 11067
rect 14105 11033 14139 11067
rect 14841 11033 14875 11067
rect 15209 11033 15243 11067
rect 4077 10965 4111 10999
rect 6929 10965 6963 10999
rect 12449 10965 12483 10999
rect 12541 10965 12575 10999
rect 13553 10965 13587 10999
rect 14749 10965 14783 10999
rect 1593 10761 1627 10795
rect 8677 10761 8711 10795
rect 10885 10761 10919 10795
rect 11529 10761 11563 10795
rect 11713 10761 11747 10795
rect 15025 10761 15059 10795
rect 8769 10693 8803 10727
rect 14657 10693 14691 10727
rect 1409 10625 1443 10659
rect 4721 10625 4755 10659
rect 4997 10625 5031 10659
rect 5181 10625 5215 10659
rect 6929 10625 6963 10659
rect 9137 10625 9171 10659
rect 9597 10625 9631 10659
rect 11667 10625 11701 10659
rect 12265 10625 12299 10659
rect 14933 10625 14967 10659
rect 1961 10557 1995 10591
rect 2237 10557 2271 10591
rect 3709 10557 3743 10591
rect 4445 10557 4479 10591
rect 4629 10557 4663 10591
rect 7205 10557 7239 10591
rect 12173 10557 12207 10591
rect 13185 10557 13219 10591
rect 15577 10557 15611 10591
rect 12081 10489 12115 10523
rect 3801 10421 3835 10455
rect 12357 10421 12391 10455
rect 2789 10217 2823 10251
rect 5549 10217 5583 10251
rect 7113 10217 7147 10251
rect 7849 10217 7883 10251
rect 12541 10217 12575 10251
rect 3433 10081 3467 10115
rect 7665 10081 7699 10115
rect 8493 10081 8527 10115
rect 9781 10081 9815 10115
rect 10057 10081 10091 10115
rect 11529 10081 11563 10115
rect 11897 10081 11931 10115
rect 14841 10081 14875 10115
rect 15117 10081 15151 10115
rect 2914 10013 2948 10047
rect 3341 10013 3375 10047
rect 8033 10013 8067 10047
rect 8217 10013 8251 10047
rect 8309 10013 8343 10047
rect 8401 10013 8435 10047
rect 8585 10013 8619 10047
rect 14105 10013 14139 10047
rect 15025 10013 15059 10047
rect 15209 10013 15243 10047
rect 15301 10013 15335 10047
rect 7021 9945 7055 9979
rect 14749 9945 14783 9979
rect 2973 9877 3007 9911
rect 4261 9673 4295 9707
rect 15117 9673 15151 9707
rect 3525 9605 3559 9639
rect 5273 9605 5307 9639
rect 11621 9605 11655 9639
rect 13645 9605 13679 9639
rect 3249 9537 3283 9571
rect 3801 9537 3835 9571
rect 3893 9537 3927 9571
rect 4202 9537 4236 9571
rect 4997 9537 5031 9571
rect 5089 9537 5123 9571
rect 5181 9537 5215 9571
rect 5457 9537 5491 9571
rect 8769 9537 8803 9571
rect 10885 9537 10919 9571
rect 11253 9537 11287 9571
rect 11805 9537 11839 9571
rect 13369 9537 13403 9571
rect 4721 9469 4755 9503
rect 4813 9469 4847 9503
rect 5549 9469 5583 9503
rect 11069 9469 11103 9503
rect 12081 9469 12115 9503
rect 4077 9333 4111 9367
rect 4629 9333 4663 9367
rect 4905 9333 4939 9367
rect 10241 9333 10275 9367
rect 11161 9333 11195 9367
rect 11989 9333 12023 9367
rect 4629 9129 4663 9163
rect 5549 9129 5583 9163
rect 8125 9129 8159 9163
rect 10057 9129 10091 9163
rect 14749 9129 14783 9163
rect 15485 9129 15519 9163
rect 8677 9061 8711 9095
rect 12265 9061 12299 9095
rect 13461 9061 13495 9095
rect 13553 9061 13587 9095
rect 2145 8993 2179 9027
rect 10885 8993 10919 9027
rect 10977 8993 11011 9027
rect 11253 8993 11287 9027
rect 11354 8993 11388 9027
rect 13093 8993 13127 9027
rect 13277 8993 13311 9027
rect 14590 8993 14624 9027
rect 1869 8925 1903 8959
rect 4077 8925 4111 8959
rect 4905 8925 4939 8959
rect 7113 8925 7147 8959
rect 7297 8925 7331 8959
rect 8033 8925 8067 8959
rect 8401 8925 8435 8959
rect 8493 8925 8527 8959
rect 9505 8925 9539 8959
rect 9873 8925 9907 8959
rect 10149 8925 10183 8959
rect 11161 8919 11195 8953
rect 11454 8925 11488 8959
rect 11621 8925 11655 8959
rect 12173 8925 12207 8959
rect 13001 8925 13035 8959
rect 14105 8925 14139 8959
rect 14841 8925 14875 8959
rect 15025 8925 15059 8959
rect 7389 8857 7423 8891
rect 12081 8857 12115 8891
rect 12449 8857 12483 8891
rect 12541 8857 12575 8891
rect 13921 8857 13955 8891
rect 14473 8857 14507 8891
rect 15577 8857 15611 8891
rect 3617 8789 3651 8823
rect 7297 8789 7331 8823
rect 8309 8789 8343 8823
rect 8953 8789 8987 8823
rect 9689 8789 9723 8823
rect 10241 8789 10275 8823
rect 12633 8789 12667 8823
rect 14381 8789 14415 8823
rect 14933 8789 14967 8823
rect 4537 8585 4571 8619
rect 9413 8585 9447 8619
rect 12173 8585 12207 8619
rect 12449 8585 12483 8619
rect 14473 8585 14507 8619
rect 8309 8517 8343 8551
rect 9137 8517 9171 8551
rect 9873 8517 9907 8551
rect 13001 8517 13035 8551
rect 15485 8517 15519 8551
rect 2789 8449 2823 8483
rect 4813 8449 4847 8483
rect 6377 8449 6411 8483
rect 9321 8449 9355 8483
rect 9505 8449 9539 8483
rect 12265 8449 12299 8483
rect 3065 8381 3099 8415
rect 4629 8381 4663 8415
rect 5089 8381 5123 8415
rect 6653 8381 6687 8415
rect 9597 8381 9631 8415
rect 11529 8381 11563 8415
rect 12725 8381 12759 8415
rect 14657 8381 14691 8415
rect 4997 8245 5031 8279
rect 8125 8245 8159 8279
rect 11345 8245 11379 8279
rect 3433 8041 3467 8075
rect 4721 8041 4755 8075
rect 8217 8041 8251 8075
rect 8677 8041 8711 8075
rect 10701 8041 10735 8075
rect 11069 7973 11103 8007
rect 13921 7973 13955 8007
rect 3617 7905 3651 7939
rect 4353 7905 4387 7939
rect 6285 7905 6319 7939
rect 6561 7905 6595 7939
rect 8953 7905 8987 7939
rect 9229 7905 9263 7939
rect 11345 7905 11379 7939
rect 12449 7905 12483 7939
rect 14841 7905 14875 7939
rect 3341 7837 3375 7871
rect 4077 7837 4111 7871
rect 4169 7837 4203 7871
rect 8401 7837 8435 7871
rect 8493 7837 8527 7871
rect 8769 7837 8803 7871
rect 10793 7837 10827 7871
rect 11161 7837 11195 7871
rect 12173 7837 12207 7871
rect 14749 7837 14783 7871
rect 6193 7769 6227 7803
rect 3617 7701 3651 7735
rect 4353 7701 4387 7735
rect 8033 7701 8067 7735
rect 14105 7701 14139 7735
rect 15485 7701 15519 7735
rect 4445 7497 4479 7531
rect 5733 7497 5767 7531
rect 8217 7497 8251 7531
rect 9689 7497 9723 7531
rect 11621 7497 11655 7531
rect 5273 7429 5307 7463
rect 9505 7429 9539 7463
rect 14473 7429 14507 7463
rect 14841 7429 14875 7463
rect 2145 7361 2179 7395
rect 4077 7361 4111 7395
rect 4353 7361 4387 7395
rect 4537 7361 4571 7395
rect 5089 7361 5123 7395
rect 5365 7361 5399 7395
rect 5825 7361 5859 7395
rect 6469 7361 6503 7395
rect 8953 7361 8987 7395
rect 9137 7361 9171 7395
rect 9597 7361 9631 7395
rect 9689 7361 9723 7395
rect 9873 7361 9907 7395
rect 11713 7361 11747 7395
rect 14749 7361 14783 7395
rect 15025 7361 15059 7395
rect 15117 7361 15151 7395
rect 15393 7361 15427 7395
rect 15485 7361 15519 7395
rect 2421 7293 2455 7327
rect 4169 7293 4203 7327
rect 5641 7293 5675 7327
rect 6745 7293 6779 7327
rect 13001 7293 13035 7327
rect 15301 7293 15335 7327
rect 5089 7225 5123 7259
rect 15577 7225 15611 7259
rect 3893 7157 3927 7191
rect 4813 7157 4847 7191
rect 6193 7157 6227 7191
rect 8401 7157 8435 7191
rect 9321 7157 9355 7191
rect 2132 6953 2166 6987
rect 4905 6953 4939 6987
rect 5641 6953 5675 6987
rect 7573 6953 7607 6987
rect 10504 6953 10538 6987
rect 11989 6953 12023 6987
rect 14105 6953 14139 6987
rect 3985 6885 4019 6919
rect 14749 6885 14783 6919
rect 1869 6817 1903 6851
rect 4813 6817 4847 6851
rect 5365 6817 5399 6851
rect 7021 6817 7055 6851
rect 7389 6817 7423 6851
rect 8033 6817 8067 6851
rect 10241 6817 10275 6851
rect 4077 6749 4111 6783
rect 4169 6749 4203 6783
rect 5089 6749 5123 6783
rect 5181 6749 5215 6783
rect 5273 6749 5307 6783
rect 5549 6749 5583 6783
rect 5641 6749 5675 6783
rect 6009 6749 6043 6783
rect 6745 6749 6779 6783
rect 7297 6749 7331 6783
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 8125 6749 8159 6783
rect 12725 6749 12759 6783
rect 14289 6749 14323 6783
rect 14565 6749 14599 6783
rect 15025 6749 15059 6783
rect 5733 6681 5767 6715
rect 5917 6681 5951 6715
rect 14749 6681 14783 6715
rect 3617 6613 3651 6647
rect 6193 6613 6227 6647
rect 12173 6613 12207 6647
rect 14473 6613 14507 6647
rect 14933 6613 14967 6647
rect 3433 6409 3467 6443
rect 5181 6409 5215 6443
rect 11529 6409 11563 6443
rect 3433 6273 3467 6307
rect 3801 6273 3835 6307
rect 4629 6273 4663 6307
rect 4905 6273 4939 6307
rect 4997 6273 5031 6307
rect 7205 6273 7239 6307
rect 7389 6273 7423 6307
rect 9597 6273 9631 6307
rect 11713 6273 11747 6307
rect 11989 6273 12023 6307
rect 12173 6273 12207 6307
rect 3249 6205 3283 6239
rect 3985 6205 4019 6239
rect 9873 6205 9907 6239
rect 11345 6205 11379 6239
rect 4537 6069 4571 6103
rect 4721 6069 4755 6103
rect 7297 6069 7331 6103
rect 10149 5865 10183 5899
rect 3157 5797 3191 5831
rect 4077 5797 4111 5831
rect 12541 5797 12575 5831
rect 6929 5729 6963 5763
rect 14105 5729 14139 5763
rect 14565 5729 14599 5763
rect 3065 5661 3099 5695
rect 3249 5661 3283 5695
rect 3341 5661 3375 5695
rect 3525 5661 3559 5695
rect 3801 5661 3835 5695
rect 6745 5661 6779 5695
rect 7113 5661 7147 5695
rect 10333 5661 10367 5695
rect 10425 5661 10459 5695
rect 12265 5661 12299 5695
rect 12357 5661 12391 5695
rect 14289 5661 14323 5695
rect 14381 5661 14415 5695
rect 14473 5661 14507 5695
rect 14657 5661 14691 5695
rect 15393 5661 15427 5695
rect 3893 5593 3927 5627
rect 4077 5593 4111 5627
rect 12541 5593 12575 5627
rect 14841 5593 14875 5627
rect 2881 5525 2915 5559
rect 6837 5525 6871 5559
rect 7021 5525 7055 5559
rect 11713 5525 11747 5559
rect 14105 5525 14139 5559
rect 3065 5321 3099 5355
rect 4445 5321 4479 5355
rect 11529 5321 11563 5355
rect 11897 5321 11931 5355
rect 15301 5321 15335 5355
rect 6101 5253 6135 5287
rect 13829 5253 13863 5287
rect 2973 5185 3007 5219
rect 3709 5185 3743 5219
rect 4721 5185 4755 5219
rect 6193 5185 6227 5219
rect 6377 5185 6411 5219
rect 6745 5185 6779 5219
rect 6929 5185 6963 5219
rect 7389 5185 7423 5219
rect 7573 5185 7607 5219
rect 7665 5185 7699 5219
rect 7757 5185 7791 5219
rect 10057 5185 10091 5219
rect 10977 5185 11011 5219
rect 11253 5185 11287 5219
rect 12541 5185 12575 5219
rect 12817 5185 12851 5219
rect 13001 5185 13035 5219
rect 13093 5185 13127 5219
rect 13553 5185 13587 5219
rect 2697 5117 2731 5151
rect 3801 5117 3835 5151
rect 7941 5147 7975 5181
rect 9873 5117 9907 5151
rect 10701 5117 10735 5151
rect 10885 5117 10919 5151
rect 11989 5117 12023 5151
rect 12081 5117 12115 5151
rect 12725 5117 12759 5151
rect 2881 5049 2915 5083
rect 6469 5049 6503 5083
rect 10793 5049 10827 5083
rect 2789 4981 2823 5015
rect 4629 4981 4663 5015
rect 7205 4981 7239 5015
rect 7849 4981 7883 5015
rect 9229 4981 9263 5015
rect 11161 4981 11195 5015
rect 12357 4981 12391 5015
rect 12817 4981 12851 5015
rect 3617 4777 3651 4811
rect 4077 4777 4111 4811
rect 4813 4777 4847 4811
rect 4997 4777 5031 4811
rect 5273 4777 5307 4811
rect 5365 4777 5399 4811
rect 10701 4777 10735 4811
rect 12541 4777 12575 4811
rect 14105 4777 14139 4811
rect 14841 4777 14875 4811
rect 8401 4709 8435 4743
rect 13645 4709 13679 4743
rect 1869 4641 1903 4675
rect 2145 4641 2179 4675
rect 5181 4641 5215 4675
rect 6561 4641 6595 4675
rect 6837 4641 6871 4675
rect 8953 4641 8987 4675
rect 9229 4641 9263 4675
rect 10977 4641 11011 4675
rect 13093 4641 13127 4675
rect 14657 4641 14691 4675
rect 3801 4573 3835 4607
rect 4077 4573 4111 4607
rect 4261 4573 4295 4607
rect 4353 4573 4387 4607
rect 4537 4573 4571 4607
rect 4905 4573 4939 4607
rect 5089 4573 5123 4607
rect 5457 4573 5491 4607
rect 6101 4573 6135 4607
rect 8401 4573 8435 4607
rect 8677 4573 8711 4607
rect 10793 4573 10827 4607
rect 11161 4573 11195 4607
rect 11529 4573 11563 4607
rect 12173 4573 12207 4607
rect 12357 4573 12391 4607
rect 12541 4573 12575 4607
rect 13277 4573 13311 4607
rect 13921 4573 13955 4607
rect 14289 4573 14323 4607
rect 14381 4573 14415 4607
rect 14473 4573 14507 4607
rect 14933 4573 14967 4607
rect 15025 4573 15059 4607
rect 4629 4437 4663 4471
rect 5549 4437 5583 4471
rect 8309 4437 8343 4471
rect 8585 4437 8619 4471
rect 11621 4437 11655 4471
rect 12725 4437 12759 4471
rect 13185 4437 13219 4471
rect 13737 4437 13771 4471
rect 14657 4437 14691 4471
rect 15669 4437 15703 4471
rect 3617 4233 3651 4267
rect 4077 4233 4111 4267
rect 6009 4233 6043 4267
rect 11253 4233 11287 4267
rect 14749 4233 14783 4267
rect 15485 4233 15519 4267
rect 11897 4165 11931 4199
rect 1869 4097 1903 4131
rect 3709 4097 3743 4131
rect 3893 4097 3927 4131
rect 4169 4097 4203 4131
rect 6377 4097 6411 4131
rect 8493 4097 8527 4131
rect 9505 4097 9539 4131
rect 11805 4097 11839 4131
rect 11989 4097 12023 4131
rect 12541 4097 12575 4131
rect 12633 4097 12667 4131
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 15025 4097 15059 4131
rect 15393 4097 15427 4131
rect 2145 4029 2179 4063
rect 3801 4029 3835 4063
rect 4261 4029 4295 4063
rect 4537 4029 4571 4063
rect 6653 4029 6687 4063
rect 9137 4029 9171 4063
rect 9781 4029 9815 4063
rect 11529 4029 11563 4063
rect 12357 4029 12391 4063
rect 13277 4029 13311 4063
rect 14841 4029 14875 4063
rect 15301 4029 15335 4063
rect 11621 3961 11655 3995
rect 12265 3961 12299 3995
rect 15209 3961 15243 3995
rect 8125 3893 8159 3927
rect 12817 3893 12851 3927
rect 4905 3689 4939 3723
rect 5733 3689 5767 3723
rect 6101 3689 6135 3723
rect 7941 3689 7975 3723
rect 9321 3689 9355 3723
rect 10228 3689 10262 3723
rect 13921 3689 13955 3723
rect 11897 3621 11931 3655
rect 15485 3621 15519 3655
rect 1869 3553 1903 3587
rect 3617 3553 3651 3587
rect 4353 3553 4387 3587
rect 4813 3553 4847 3587
rect 5273 3553 5307 3587
rect 6193 3553 6227 3587
rect 6469 3553 6503 3587
rect 8677 3553 8711 3587
rect 9413 3553 9447 3587
rect 9965 3553 9999 3587
rect 12173 3553 12207 3587
rect 4997 3485 5031 3519
rect 5089 3485 5123 3519
rect 5181 3485 5215 3519
rect 5365 3485 5399 3519
rect 5641 3485 5675 3519
rect 5917 3485 5951 3519
rect 8217 3485 8251 3519
rect 8309 3485 8343 3519
rect 8493 3485 8527 3519
rect 9137 3485 9171 3519
rect 9229 3485 9263 3519
rect 11989 3485 12023 3519
rect 14749 3485 14783 3519
rect 14933 3485 14967 3519
rect 2145 3417 2179 3451
rect 12449 3417 12483 3451
rect 14105 3417 14139 3451
rect 3801 3349 3835 3383
rect 11713 3349 11747 3383
rect 2881 3145 2915 3179
rect 6469 3145 6503 3179
rect 10241 3145 10275 3179
rect 10977 3145 11011 3179
rect 13001 3145 13035 3179
rect 13369 3077 13403 3111
rect 14933 3077 14967 3111
rect 3065 3009 3099 3043
rect 3249 3009 3283 3043
rect 3525 3009 3559 3043
rect 7021 3009 7055 3043
rect 7205 3009 7239 3043
rect 7297 3009 7331 3043
rect 7573 3009 7607 3043
rect 7849 3009 7883 3043
rect 7941 3009 7975 3043
rect 10425 3009 10459 3043
rect 10517 3009 10551 3043
rect 10793 3009 10827 3043
rect 11069 3009 11103 3043
rect 12357 3009 12391 3043
rect 13093 3009 13127 3043
rect 15117 3009 15151 3043
rect 15301 3009 15335 3043
rect 3341 2941 3375 2975
rect 15393 2941 15427 2975
rect 3157 2873 3191 2907
rect 10701 2873 10735 2907
rect 14841 2805 14875 2839
rect 14657 2601 14691 2635
rect 1685 2533 1719 2567
rect 14749 2533 14783 2567
rect 15117 2465 15151 2499
rect 9873 2397 9907 2431
rect 13093 2397 13127 2431
rect 1501 2329 1535 2363
rect 9965 2261 9999 2295
rect 13185 2261 13219 2295
<< metal1 >>
rect 1104 16890 16008 16912
rect 1104 16838 2813 16890
rect 2865 16838 2877 16890
rect 2929 16838 2941 16890
rect 2993 16838 3005 16890
rect 3057 16838 3069 16890
rect 3121 16838 6539 16890
rect 6591 16838 6603 16890
rect 6655 16838 6667 16890
rect 6719 16838 6731 16890
rect 6783 16838 6795 16890
rect 6847 16838 10265 16890
rect 10317 16838 10329 16890
rect 10381 16838 10393 16890
rect 10445 16838 10457 16890
rect 10509 16838 10521 16890
rect 10573 16838 13991 16890
rect 14043 16838 14055 16890
rect 14107 16838 14119 16890
rect 14171 16838 14183 16890
rect 14235 16838 14247 16890
rect 14299 16838 16008 16890
rect 1104 16816 16008 16838
rect 7392 16680 8156 16708
rect 7392 16649 7420 16680
rect 8128 16652 8156 16680
rect 7377 16643 7435 16649
rect 7377 16609 7389 16643
rect 7423 16609 7435 16643
rect 7377 16603 7435 16609
rect 7469 16643 7527 16649
rect 7469 16609 7481 16643
rect 7515 16640 7527 16643
rect 7837 16643 7895 16649
rect 7837 16640 7849 16643
rect 7515 16612 7849 16640
rect 7515 16609 7527 16612
rect 7469 16603 7527 16609
rect 7837 16609 7849 16612
rect 7883 16609 7895 16643
rect 7837 16603 7895 16609
rect 8110 16600 8116 16652
rect 8168 16600 8174 16652
rect 8386 16600 8392 16652
rect 8444 16600 8450 16652
rect 11422 16600 11428 16652
rect 11480 16640 11486 16652
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11480 16612 11897 16640
rect 11480 16600 11486 16612
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 12069 16643 12127 16649
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 12894 16640 12900 16652
rect 12115 16612 12900 16640
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 12894 16600 12900 16612
rect 12952 16600 12958 16652
rect 5350 16532 5356 16584
rect 5408 16532 5414 16584
rect 7561 16575 7619 16581
rect 7561 16541 7573 16575
rect 7607 16541 7619 16575
rect 7561 16535 7619 16541
rect 7576 16504 7604 16535
rect 7650 16532 7656 16584
rect 7708 16532 7714 16584
rect 11330 16532 11336 16584
rect 11388 16572 11394 16584
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 11388 16544 11805 16572
rect 11388 16532 11394 16544
rect 11793 16541 11805 16544
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 11977 16575 12035 16581
rect 11977 16541 11989 16575
rect 12023 16572 12035 16575
rect 12342 16572 12348 16584
rect 12023 16544 12348 16572
rect 12023 16541 12035 16544
rect 11977 16535 12035 16541
rect 12342 16532 12348 16544
rect 12400 16532 12406 16584
rect 7576 16476 7696 16504
rect 4338 16396 4344 16448
rect 4396 16436 4402 16448
rect 4801 16439 4859 16445
rect 4801 16436 4813 16439
rect 4396 16408 4813 16436
rect 4396 16396 4402 16408
rect 4801 16405 4813 16408
rect 4847 16405 4859 16439
rect 4801 16399 4859 16405
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 7193 16439 7251 16445
rect 7193 16436 7205 16439
rect 7156 16408 7205 16436
rect 7156 16396 7162 16408
rect 7193 16405 7205 16408
rect 7239 16405 7251 16439
rect 7668 16436 7696 16476
rect 9122 16436 9128 16448
rect 7668 16408 9128 16436
rect 7193 16399 7251 16405
rect 9122 16396 9128 16408
rect 9180 16396 9186 16448
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 11609 16439 11667 16445
rect 11609 16436 11621 16439
rect 10836 16408 11621 16436
rect 10836 16396 10842 16408
rect 11609 16405 11621 16408
rect 11655 16405 11667 16439
rect 11609 16399 11667 16405
rect 1104 16346 16008 16368
rect 1104 16294 3473 16346
rect 3525 16294 3537 16346
rect 3589 16294 3601 16346
rect 3653 16294 3665 16346
rect 3717 16294 3729 16346
rect 3781 16294 7199 16346
rect 7251 16294 7263 16346
rect 7315 16294 7327 16346
rect 7379 16294 7391 16346
rect 7443 16294 7455 16346
rect 7507 16294 10925 16346
rect 10977 16294 10989 16346
rect 11041 16294 11053 16346
rect 11105 16294 11117 16346
rect 11169 16294 11181 16346
rect 11233 16294 14651 16346
rect 14703 16294 14715 16346
rect 14767 16294 14779 16346
rect 14831 16294 14843 16346
rect 14895 16294 14907 16346
rect 14959 16294 16008 16346
rect 1104 16272 16008 16294
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5350 16232 5356 16244
rect 5040 16204 5356 16232
rect 5040 16192 5046 16204
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 7098 16192 7104 16244
rect 7156 16192 7162 16244
rect 9122 16192 9128 16244
rect 9180 16232 9186 16244
rect 9677 16235 9735 16241
rect 9677 16232 9689 16235
rect 9180 16204 9689 16232
rect 9180 16192 9186 16204
rect 9677 16201 9689 16204
rect 9723 16232 9735 16235
rect 11422 16232 11428 16244
rect 9723 16204 11428 16232
rect 9723 16201 9735 16204
rect 9677 16195 9735 16201
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 5994 16096 6000 16108
rect 4646 16068 6000 16096
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 7116 16105 7144 16192
rect 10134 16164 10140 16176
rect 9430 16136 10140 16164
rect 10134 16124 10140 16136
rect 10192 16124 10198 16176
rect 10778 16124 10784 16176
rect 10836 16164 10842 16176
rect 11241 16167 11299 16173
rect 10836 16136 10916 16164
rect 10836 16124 10842 16136
rect 10888 16105 10916 16136
rect 11241 16133 11253 16167
rect 11287 16164 11299 16167
rect 12345 16167 12403 16173
rect 12345 16164 12357 16167
rect 11287 16136 12357 16164
rect 11287 16133 11299 16136
rect 11241 16127 11299 16133
rect 12345 16133 12357 16136
rect 12391 16164 12403 16167
rect 12434 16164 12440 16176
rect 12391 16136 12440 16164
rect 12391 16133 12403 16136
rect 12345 16127 12403 16133
rect 12434 16124 12440 16136
rect 12492 16124 12498 16176
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 10873 16099 10931 16105
rect 10873 16065 10885 16099
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 11333 16100 11391 16105
rect 11333 16099 11468 16100
rect 11333 16065 11345 16099
rect 11379 16096 11468 16099
rect 11379 16072 12388 16096
rect 11379 16065 11391 16072
rect 11440 16068 12388 16072
rect 11333 16059 11391 16065
rect 12360 16040 12388 16068
rect 12894 16056 12900 16108
rect 12952 16056 12958 16108
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 15997 3295 16031
rect 3237 15991 3295 15997
rect 3513 16031 3571 16037
rect 3513 15997 3525 16031
rect 3559 16028 3571 16031
rect 3878 16028 3884 16040
rect 3559 16000 3884 16028
rect 3559 15997 3571 16000
rect 3513 15991 3571 15997
rect 3252 15892 3280 15991
rect 3878 15988 3884 16000
rect 3936 15988 3942 16040
rect 5534 15988 5540 16040
rect 5592 16028 5598 16040
rect 5629 16031 5687 16037
rect 5629 16028 5641 16031
rect 5592 16000 5641 16028
rect 5592 15988 5598 16000
rect 5629 15997 5641 16000
rect 5675 15997 5687 16031
rect 5629 15991 5687 15997
rect 7926 15988 7932 16040
rect 7984 15988 7990 16040
rect 8202 15988 8208 16040
rect 8260 15988 8266 16040
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 16028 11115 16031
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 11103 16000 11529 16028
rect 11103 15997 11115 16000
rect 11057 15991 11115 15997
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 11517 15991 11575 15997
rect 12342 15988 12348 16040
rect 12400 15988 12406 16040
rect 4614 15892 4620 15904
rect 3252 15864 4620 15892
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 5074 15852 5080 15904
rect 5132 15852 5138 15904
rect 7653 15895 7711 15901
rect 7653 15861 7665 15895
rect 7699 15892 7711 15895
rect 7834 15892 7840 15904
rect 7699 15864 7840 15892
rect 7699 15861 7711 15864
rect 7653 15855 7711 15861
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 12158 15852 12164 15904
rect 12216 15852 12222 15904
rect 1104 15802 16008 15824
rect 1104 15750 2813 15802
rect 2865 15750 2877 15802
rect 2929 15750 2941 15802
rect 2993 15750 3005 15802
rect 3057 15750 3069 15802
rect 3121 15750 6539 15802
rect 6591 15750 6603 15802
rect 6655 15750 6667 15802
rect 6719 15750 6731 15802
rect 6783 15750 6795 15802
rect 6847 15750 10265 15802
rect 10317 15750 10329 15802
rect 10381 15750 10393 15802
rect 10445 15750 10457 15802
rect 10509 15750 10521 15802
rect 10573 15750 13991 15802
rect 14043 15750 14055 15802
rect 14107 15750 14119 15802
rect 14171 15750 14183 15802
rect 14235 15750 14247 15802
rect 14299 15750 16008 15802
rect 1104 15728 16008 15750
rect 4880 15691 4938 15697
rect 4880 15657 4892 15691
rect 4926 15688 4938 15691
rect 5074 15688 5080 15700
rect 4926 15660 5080 15688
rect 4926 15657 4938 15660
rect 4880 15651 4938 15657
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 7941 15691 7999 15697
rect 7941 15688 7953 15691
rect 7892 15660 7953 15688
rect 7892 15648 7898 15660
rect 7941 15657 7953 15660
rect 7987 15657 7999 15691
rect 7941 15651 7999 15657
rect 8202 15648 8208 15700
rect 8260 15688 8266 15700
rect 8297 15691 8355 15697
rect 8297 15688 8309 15691
rect 8260 15660 8309 15688
rect 8260 15648 8266 15660
rect 8297 15657 8309 15660
rect 8343 15657 8355 15691
rect 8297 15651 8355 15657
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10192 15660 12848 15688
rect 10192 15648 10198 15660
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15552 1915 15555
rect 4614 15552 4620 15564
rect 1903 15524 4620 15552
rect 1903 15521 1915 15524
rect 1857 15515 1915 15521
rect 4614 15512 4620 15524
rect 4672 15552 4678 15564
rect 7926 15552 7932 15564
rect 4672 15524 7932 15552
rect 4672 15512 4678 15524
rect 6932 15496 6960 15524
rect 7926 15512 7932 15524
rect 7984 15552 7990 15564
rect 8205 15555 8263 15561
rect 8205 15552 8217 15555
rect 7984 15524 8217 15552
rect 7984 15512 7990 15524
rect 8205 15521 8217 15524
rect 8251 15521 8263 15555
rect 10137 15555 10195 15561
rect 8205 15515 8263 15521
rect 9784 15524 9996 15552
rect 9784 15496 9812 15524
rect 3789 15487 3847 15493
rect 3789 15484 3801 15487
rect 3620 15456 3801 15484
rect 2133 15419 2191 15425
rect 2133 15385 2145 15419
rect 2179 15385 2191 15419
rect 2133 15379 2191 15385
rect 2148 15348 2176 15379
rect 3142 15376 3148 15428
rect 3200 15376 3206 15428
rect 2774 15348 2780 15360
rect 2148 15320 2780 15348
rect 2774 15308 2780 15320
rect 2832 15308 2838 15360
rect 3620 15357 3648 15456
rect 3789 15453 3801 15456
rect 3835 15453 3847 15487
rect 3789 15447 3847 15453
rect 5994 15444 6000 15496
rect 6052 15484 6058 15496
rect 6052 15456 6854 15484
rect 6052 15444 6058 15456
rect 6914 15444 6920 15496
rect 6972 15444 6978 15496
rect 8478 15444 8484 15496
rect 8536 15444 8542 15496
rect 9766 15444 9772 15496
rect 9824 15444 9830 15496
rect 9858 15444 9864 15496
rect 9916 15444 9922 15496
rect 9968 15493 9996 15524
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 11422 15552 11428 15564
rect 10183 15524 11428 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 11793 15555 11851 15561
rect 11793 15521 11805 15555
rect 11839 15552 11851 15555
rect 12158 15552 12164 15564
rect 11839 15524 12164 15552
rect 11839 15521 11851 15524
rect 11793 15515 11851 15521
rect 12158 15512 12164 15524
rect 12216 15512 12222 15564
rect 9953 15487 10011 15493
rect 9953 15453 9965 15487
rect 9999 15453 10011 15487
rect 9953 15447 10011 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15484 10287 15487
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10275 15456 10701 15484
rect 10275 15453 10287 15456
rect 10229 15447 10287 15453
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 11330 15444 11336 15496
rect 11388 15444 11394 15496
rect 11517 15487 11575 15493
rect 11517 15453 11529 15487
rect 11563 15453 11575 15487
rect 12820 15484 12848 15660
rect 12894 15648 12900 15700
rect 12952 15688 12958 15700
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 12952 15660 13277 15688
rect 12952 15648 12958 15660
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 12894 15484 12900 15496
rect 12820 15456 12900 15484
rect 11517 15447 11575 15453
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15317 3663 15351
rect 3605 15311 3663 15317
rect 4246 15308 4252 15360
rect 4304 15348 4310 15360
rect 4433 15351 4491 15357
rect 4433 15348 4445 15351
rect 4304 15320 4445 15348
rect 4304 15308 4310 15320
rect 4433 15317 4445 15320
rect 4479 15317 4491 15351
rect 4433 15311 4491 15317
rect 5626 15308 5632 15360
rect 5684 15348 5690 15360
rect 6362 15348 6368 15360
rect 5684 15320 6368 15348
rect 5684 15308 5690 15320
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 6457 15351 6515 15357
rect 6457 15317 6469 15351
rect 6503 15348 6515 15351
rect 6546 15348 6552 15360
rect 6503 15320 6552 15348
rect 6503 15317 6515 15320
rect 6457 15311 6515 15317
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 9674 15308 9680 15360
rect 9732 15308 9738 15360
rect 11532 15348 11560 15447
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 13280 15456 13553 15484
rect 13280 15360 13308 15456
rect 13541 15453 13553 15456
rect 13587 15453 13599 15487
rect 13541 15447 13599 15453
rect 11974 15348 11980 15360
rect 11532 15320 11980 15348
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 13262 15308 13268 15360
rect 13320 15308 13326 15360
rect 13446 15308 13452 15360
rect 13504 15308 13510 15360
rect 1104 15258 16008 15280
rect 1104 15206 3473 15258
rect 3525 15206 3537 15258
rect 3589 15206 3601 15258
rect 3653 15206 3665 15258
rect 3717 15206 3729 15258
rect 3781 15206 7199 15258
rect 7251 15206 7263 15258
rect 7315 15206 7327 15258
rect 7379 15206 7391 15258
rect 7443 15206 7455 15258
rect 7507 15206 10925 15258
rect 10977 15206 10989 15258
rect 11041 15206 11053 15258
rect 11105 15206 11117 15258
rect 11169 15206 11181 15258
rect 11233 15206 14651 15258
rect 14703 15206 14715 15258
rect 14767 15206 14779 15258
rect 14831 15206 14843 15258
rect 14895 15206 14907 15258
rect 14959 15206 16008 15258
rect 1104 15184 16008 15206
rect 3878 15104 3884 15156
rect 3936 15104 3942 15156
rect 5000 15116 6316 15144
rect 5000 15088 5028 15116
rect 4614 15076 4620 15088
rect 3252 15048 4292 15076
rect 3252 15017 3280 15048
rect 4264 15020 4292 15048
rect 4448 15048 4620 15076
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 3237 15011 3295 15017
rect 3237 15008 3249 15011
rect 3007 14980 3249 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 3237 14977 3249 14980
rect 3283 14977 3295 15011
rect 3237 14971 3295 14977
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 3970 15008 3976 15020
rect 3467 14980 3976 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4065 15011 4123 15017
rect 4065 14977 4077 15011
rect 4111 14977 4123 15011
rect 4065 14971 4123 14977
rect 2685 14943 2743 14949
rect 2685 14909 2697 14943
rect 2731 14940 2743 14943
rect 3329 14943 3387 14949
rect 3329 14940 3341 14943
rect 2731 14912 3341 14940
rect 2731 14909 2743 14912
rect 2685 14903 2743 14909
rect 3329 14909 3341 14912
rect 3375 14909 3387 14943
rect 3329 14903 3387 14909
rect 2774 14832 2780 14884
rect 2832 14832 2838 14884
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 2869 14807 2927 14813
rect 2869 14804 2881 14807
rect 2740 14776 2881 14804
rect 2740 14764 2746 14776
rect 2869 14773 2881 14776
rect 2915 14773 2927 14807
rect 4080 14804 4108 14971
rect 4246 14968 4252 15020
rect 4304 14968 4310 15020
rect 4448 15017 4476 15048
rect 4614 15036 4620 15048
rect 4672 15036 4678 15088
rect 4982 15036 4988 15088
rect 5040 15036 5046 15088
rect 6288 15076 6316 15116
rect 6362 15104 6368 15156
rect 6420 15144 6426 15156
rect 6917 15147 6975 15153
rect 6917 15144 6929 15147
rect 6420 15116 6929 15144
rect 6420 15104 6426 15116
rect 6917 15113 6929 15116
rect 6963 15113 6975 15147
rect 6917 15107 6975 15113
rect 7193 15147 7251 15153
rect 7193 15113 7205 15147
rect 7239 15144 7251 15147
rect 7650 15144 7656 15156
rect 7239 15116 7656 15144
rect 7239 15113 7251 15116
rect 7193 15107 7251 15113
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 8297 15147 8355 15153
rect 8297 15113 8309 15147
rect 8343 15144 8355 15147
rect 8386 15144 8392 15156
rect 8343 15116 8392 15144
rect 8343 15113 8355 15116
rect 8297 15107 8355 15113
rect 7034 15079 7092 15085
rect 7034 15076 7046 15079
rect 6288 15048 7046 15076
rect 7034 15045 7046 15048
rect 7080 15076 7092 15079
rect 7374 15076 7380 15088
rect 7080 15048 7380 15076
rect 7080 15045 7092 15048
rect 7034 15039 7092 15045
rect 7374 15036 7380 15048
rect 7432 15036 7438 15088
rect 4433 15011 4491 15017
rect 4433 14977 4445 15011
rect 4479 14977 4491 15011
rect 5994 15008 6000 15020
rect 5842 14980 6000 15008
rect 4433 14971 4491 14977
rect 5994 14968 6000 14980
rect 6052 14968 6058 15020
rect 6546 14968 6552 15020
rect 6604 15008 6610 15020
rect 8312 15008 8340 15107
rect 8386 15104 8392 15116
rect 8444 15104 8450 15156
rect 8478 15104 8484 15156
rect 8536 15144 8542 15156
rect 8757 15147 8815 15153
rect 8757 15144 8769 15147
rect 8536 15116 8769 15144
rect 8536 15104 8542 15116
rect 8757 15113 8769 15116
rect 8803 15113 8815 15147
rect 8757 15107 8815 15113
rect 9122 15104 9128 15156
rect 9180 15104 9186 15156
rect 9217 15147 9275 15153
rect 9217 15113 9229 15147
rect 9263 15144 9275 15147
rect 9263 15116 9812 15144
rect 9263 15113 9275 15116
rect 9217 15107 9275 15113
rect 6604 14980 8340 15008
rect 6604 14968 6610 14980
rect 8386 14968 8392 15020
rect 8444 14968 8450 15020
rect 9140 15017 9168 15104
rect 9125 15011 9183 15017
rect 9125 14977 9137 15011
rect 9171 14977 9183 15011
rect 9125 14971 9183 14977
rect 4338 14900 4344 14952
rect 4396 14900 4402 14952
rect 4706 14900 4712 14952
rect 4764 14900 4770 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6104 14912 6837 14940
rect 5258 14804 5264 14816
rect 4080 14776 5264 14804
rect 2869 14767 2927 14773
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 6104 14804 6132 14912
rect 6825 14909 6837 14912
rect 6871 14940 6883 14943
rect 7466 14940 7472 14952
rect 6871 14912 7472 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 7466 14900 7472 14912
rect 7524 14900 7530 14952
rect 7837 14943 7895 14949
rect 7837 14909 7849 14943
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 8205 14943 8263 14949
rect 8205 14909 8217 14943
rect 8251 14940 8263 14943
rect 8251 14912 8340 14940
rect 8251 14909 8263 14912
rect 8205 14903 8263 14909
rect 7852 14872 7880 14903
rect 6196 14844 7880 14872
rect 8312 14872 8340 14912
rect 9232 14872 9260 15107
rect 9784 15088 9812 15116
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 14458 15144 14464 15156
rect 12952 15116 13584 15144
rect 12952 15104 12958 15116
rect 9674 15036 9680 15088
rect 9732 15036 9738 15088
rect 9766 15036 9772 15088
rect 9824 15036 9830 15088
rect 10134 15036 10140 15088
rect 10192 15036 10198 15088
rect 12710 15036 12716 15088
rect 12768 15036 12774 15088
rect 13556 15076 13584 15116
rect 14016 15116 14464 15144
rect 14016 15076 14044 15116
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 13556 15048 14122 15076
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14940 9459 14943
rect 11974 14940 11980 14952
rect 9447 14912 9536 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 8312 14844 9260 14872
rect 6196 14816 6224 14844
rect 9508 14816 9536 14912
rect 10704 14912 11980 14940
rect 5500 14776 6132 14804
rect 5500 14764 5506 14776
rect 6178 14764 6184 14816
rect 6236 14764 6242 14816
rect 7282 14764 7288 14816
rect 7340 14764 7346 14816
rect 9490 14764 9496 14816
rect 9548 14804 9554 14816
rect 10704 14804 10732 14912
rect 11974 14900 11980 14912
rect 12032 14900 12038 14952
rect 12250 14900 12256 14952
rect 12308 14900 12314 14952
rect 15286 14900 15292 14952
rect 15344 14900 15350 14952
rect 15562 14900 15568 14952
rect 15620 14900 15626 14952
rect 9548 14776 10732 14804
rect 11149 14807 11207 14813
rect 9548 14764 9554 14776
rect 11149 14773 11161 14807
rect 11195 14804 11207 14807
rect 11330 14804 11336 14816
rect 11195 14776 11336 14804
rect 11195 14773 11207 14776
rect 11149 14767 11207 14773
rect 11330 14764 11336 14776
rect 11388 14804 11394 14816
rect 11514 14804 11520 14816
rect 11388 14776 11520 14804
rect 11388 14764 11394 14776
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 13725 14807 13783 14813
rect 13725 14804 13737 14807
rect 13320 14776 13737 14804
rect 13320 14764 13326 14776
rect 13725 14773 13737 14776
rect 13771 14773 13783 14807
rect 13725 14767 13783 14773
rect 13814 14764 13820 14816
rect 13872 14764 13878 14816
rect 1104 14714 16008 14736
rect 1104 14662 2813 14714
rect 2865 14662 2877 14714
rect 2929 14662 2941 14714
rect 2993 14662 3005 14714
rect 3057 14662 3069 14714
rect 3121 14662 6539 14714
rect 6591 14662 6603 14714
rect 6655 14662 6667 14714
rect 6719 14662 6731 14714
rect 6783 14662 6795 14714
rect 6847 14662 10265 14714
rect 10317 14662 10329 14714
rect 10381 14662 10393 14714
rect 10445 14662 10457 14714
rect 10509 14662 10521 14714
rect 10573 14662 13991 14714
rect 14043 14662 14055 14714
rect 14107 14662 14119 14714
rect 14171 14662 14183 14714
rect 14235 14662 14247 14714
rect 14299 14662 16008 14714
rect 1104 14640 16008 14662
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 4801 14603 4859 14609
rect 4801 14600 4813 14603
rect 4764 14572 4813 14600
rect 4764 14560 4770 14572
rect 4801 14569 4813 14572
rect 4847 14569 4859 14603
rect 4801 14563 4859 14569
rect 5445 14603 5503 14609
rect 5445 14569 5457 14603
rect 5491 14600 5503 14603
rect 7282 14600 7288 14612
rect 5491 14572 7288 14600
rect 5491 14569 5503 14572
rect 5445 14563 5503 14569
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 8297 14603 8355 14609
rect 8297 14600 8309 14603
rect 7524 14572 8309 14600
rect 7524 14560 7530 14572
rect 5077 14535 5135 14541
rect 5077 14501 5089 14535
rect 5123 14532 5135 14535
rect 5534 14532 5540 14544
rect 5123 14504 5540 14532
rect 5123 14501 5135 14504
rect 5077 14495 5135 14501
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 5629 14535 5687 14541
rect 5629 14501 5641 14535
rect 5675 14501 5687 14535
rect 5629 14495 5687 14501
rect 5644 14464 5672 14495
rect 6178 14492 6184 14544
rect 6236 14532 6242 14544
rect 6236 14504 7052 14532
rect 6236 14492 6242 14504
rect 7024 14473 7052 14504
rect 7374 14492 7380 14544
rect 7432 14532 7438 14544
rect 7432 14504 8064 14532
rect 7432 14492 7438 14504
rect 5000 14436 5672 14464
rect 6273 14467 6331 14473
rect 5000 14405 5028 14436
rect 6273 14433 6285 14467
rect 6319 14464 6331 14467
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 6319 14436 6469 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14433 7067 14467
rect 7745 14467 7803 14473
rect 7745 14464 7757 14467
rect 7009 14427 7067 14433
rect 7116 14436 7757 14464
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14365 5043 14399
rect 4985 14359 5043 14365
rect 5258 14356 5264 14408
rect 5316 14356 5322 14408
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 7116 14396 7144 14436
rect 7745 14433 7757 14436
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 5592 14368 7144 14396
rect 7285 14399 7343 14405
rect 5592 14356 5598 14368
rect 7285 14365 7297 14399
rect 7331 14396 7343 14399
rect 7374 14396 7380 14408
rect 7331 14368 7380 14396
rect 7331 14365 7343 14368
rect 7285 14359 7343 14365
rect 7374 14356 7380 14368
rect 7432 14356 7438 14408
rect 7760 14396 7788 14427
rect 7837 14399 7895 14405
rect 7837 14396 7849 14399
rect 7760 14368 7849 14396
rect 7837 14365 7849 14368
rect 7883 14365 7895 14399
rect 7837 14359 7895 14365
rect 5276 14260 5304 14356
rect 8036 14337 8064 14504
rect 8128 14405 8156 14572
rect 8297 14569 8309 14572
rect 8343 14569 8355 14603
rect 8297 14563 8355 14569
rect 9122 14560 9128 14612
rect 9180 14560 9186 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10042 14600 10048 14612
rect 9916 14572 10048 14600
rect 9916 14560 9922 14572
rect 10042 14560 10048 14572
rect 10100 14600 10106 14612
rect 11701 14603 11759 14609
rect 11701 14600 11713 14603
rect 10100 14572 11713 14600
rect 10100 14560 10106 14572
rect 11701 14569 11713 14572
rect 11747 14569 11759 14603
rect 11701 14563 11759 14569
rect 12250 14560 12256 14612
rect 12308 14560 12314 14612
rect 14737 14603 14795 14609
rect 14737 14569 14749 14603
rect 14783 14600 14795 14603
rect 15286 14600 15292 14612
rect 14783 14572 15292 14600
rect 14783 14569 14795 14572
rect 14737 14563 14795 14569
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 9140 14532 9168 14560
rect 8404 14504 9168 14532
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14365 8171 14399
rect 8113 14359 8171 14365
rect 8202 14356 8208 14408
rect 8260 14356 8266 14408
rect 8404 14405 8432 14504
rect 12986 14492 12992 14544
rect 13044 14532 13050 14544
rect 13725 14535 13783 14541
rect 13725 14532 13737 14535
rect 13044 14504 13737 14532
rect 13044 14492 13050 14504
rect 13725 14501 13737 14504
rect 13771 14532 13783 14535
rect 13771 14504 14504 14532
rect 13771 14501 13783 14504
rect 13725 14495 13783 14501
rect 8846 14424 8852 14476
rect 8904 14464 8910 14476
rect 9125 14467 9183 14473
rect 9125 14464 9137 14467
rect 8904 14436 9137 14464
rect 8904 14424 8910 14436
rect 9125 14433 9137 14436
rect 9171 14464 9183 14467
rect 9490 14464 9496 14476
rect 9171 14436 9496 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 12161 14467 12219 14473
rect 9824 14436 11008 14464
rect 9824 14424 9830 14436
rect 10980 14405 11008 14436
rect 12161 14433 12173 14467
rect 12207 14464 12219 14467
rect 13814 14464 13820 14476
rect 12207 14436 13820 14464
rect 12207 14433 12219 14436
rect 12161 14427 12219 14433
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 11609 14399 11667 14405
rect 11609 14396 11621 14399
rect 11195 14368 11621 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11609 14365 11621 14368
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 11977 14399 12035 14405
rect 11977 14365 11989 14399
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 8021 14331 8079 14337
rect 8021 14297 8033 14331
rect 8067 14297 8079 14331
rect 8021 14291 8079 14297
rect 5718 14260 5724 14272
rect 5276 14232 5724 14260
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 5902 14220 5908 14272
rect 5960 14260 5966 14272
rect 5997 14263 6055 14269
rect 5997 14260 6009 14263
rect 5960 14232 6009 14260
rect 5960 14220 5966 14232
rect 5997 14229 6009 14232
rect 6043 14229 6055 14263
rect 5997 14223 6055 14229
rect 6089 14263 6147 14269
rect 6089 14229 6101 14263
rect 6135 14260 6147 14263
rect 7006 14260 7012 14272
rect 6135 14232 7012 14260
rect 6135 14229 6147 14232
rect 6089 14223 6147 14229
rect 7006 14220 7012 14232
rect 7064 14260 7070 14272
rect 7285 14263 7343 14269
rect 7285 14260 7297 14263
rect 7064 14232 7297 14260
rect 7064 14220 7070 14232
rect 7285 14229 7297 14232
rect 7331 14229 7343 14263
rect 7285 14223 7343 14229
rect 7926 14220 7932 14272
rect 7984 14220 7990 14272
rect 8220 14260 8248 14356
rect 9398 14288 9404 14340
rect 9456 14288 9462 14340
rect 10134 14288 10140 14340
rect 10192 14288 10198 14340
rect 11514 14288 11520 14340
rect 11572 14328 11578 14340
rect 11624 14328 11652 14359
rect 11572 14300 11652 14328
rect 11992 14328 12020 14359
rect 12434 14356 12440 14408
rect 12492 14356 12498 14408
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12544 14328 12572 14359
rect 12986 14356 12992 14408
rect 13044 14396 13050 14408
rect 13081 14399 13139 14405
rect 13081 14396 13093 14399
rect 13044 14368 13093 14396
rect 13044 14356 13050 14368
rect 13081 14365 13093 14368
rect 13127 14365 13139 14399
rect 13081 14359 13139 14365
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13228 14368 13277 14396
rect 13228 14356 13234 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 13354 14356 13360 14408
rect 13412 14356 13418 14408
rect 13556 14405 13584 14436
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 14476 14405 14504 14504
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14433 14611 14467
rect 14553 14427 14611 14433
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13633 14399 13691 14405
rect 13633 14396 13645 14399
rect 13587 14368 13645 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 13633 14365 13645 14368
rect 13679 14365 13691 14399
rect 13633 14359 13691 14365
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 13372 14328 13400 14356
rect 11992 14300 13400 14328
rect 13449 14331 13507 14337
rect 11572 14288 11578 14300
rect 13449 14297 13461 14331
rect 13495 14328 13507 14331
rect 14093 14331 14151 14337
rect 14093 14328 14105 14331
rect 13495 14300 14105 14328
rect 13495 14297 13507 14300
rect 13449 14291 13507 14297
rect 13648 14272 13676 14300
rect 14093 14297 14105 14300
rect 14139 14297 14151 14331
rect 14093 14291 14151 14297
rect 10042 14260 10048 14272
rect 8220 14232 10048 14260
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 10873 14263 10931 14269
rect 10873 14260 10885 14263
rect 10744 14232 10885 14260
rect 10744 14220 10750 14232
rect 10873 14229 10885 14232
rect 10919 14229 10931 14263
rect 10873 14223 10931 14229
rect 11057 14263 11115 14269
rect 11057 14229 11069 14263
rect 11103 14260 11115 14263
rect 11330 14260 11336 14272
rect 11103 14232 11336 14260
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 12342 14220 12348 14272
rect 12400 14260 12406 14272
rect 12897 14263 12955 14269
rect 12897 14260 12909 14263
rect 12400 14232 12909 14260
rect 12400 14220 12406 14232
rect 12897 14229 12909 14232
rect 12943 14260 12955 14263
rect 13081 14263 13139 14269
rect 13081 14260 13093 14263
rect 12943 14232 13093 14260
rect 12943 14229 12955 14232
rect 12897 14223 12955 14229
rect 13081 14229 13093 14232
rect 13127 14229 13139 14263
rect 13081 14223 13139 14229
rect 13630 14220 13636 14272
rect 13688 14220 13694 14272
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 14568 14260 14596 14427
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15381 14399 15439 14405
rect 15381 14396 15393 14399
rect 15068 14368 15393 14396
rect 15068 14356 15074 14368
rect 15381 14365 15393 14368
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 14829 14263 14887 14269
rect 14829 14260 14841 14263
rect 13964 14232 14841 14260
rect 13964 14220 13970 14232
rect 14829 14229 14841 14232
rect 14875 14229 14887 14263
rect 14829 14223 14887 14229
rect 1104 14170 16008 14192
rect 1104 14118 3473 14170
rect 3525 14118 3537 14170
rect 3589 14118 3601 14170
rect 3653 14118 3665 14170
rect 3717 14118 3729 14170
rect 3781 14118 7199 14170
rect 7251 14118 7263 14170
rect 7315 14118 7327 14170
rect 7379 14118 7391 14170
rect 7443 14118 7455 14170
rect 7507 14118 10925 14170
rect 10977 14118 10989 14170
rect 11041 14118 11053 14170
rect 11105 14118 11117 14170
rect 11169 14118 11181 14170
rect 11233 14118 14651 14170
rect 14703 14118 14715 14170
rect 14767 14118 14779 14170
rect 14831 14118 14843 14170
rect 14895 14118 14907 14170
rect 14959 14118 16008 14170
rect 1104 14096 16008 14118
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 4798 14056 4804 14068
rect 4212 14028 4804 14056
rect 4212 14016 4218 14028
rect 4798 14016 4804 14028
rect 4856 14056 4862 14068
rect 5353 14059 5411 14065
rect 5353 14056 5365 14059
rect 4856 14028 5365 14056
rect 4856 14016 4862 14028
rect 5353 14025 5365 14028
rect 5399 14025 5411 14059
rect 5353 14019 5411 14025
rect 5442 14016 5448 14068
rect 5500 14016 5506 14068
rect 5718 14016 5724 14068
rect 5776 14056 5782 14068
rect 7926 14056 7932 14068
rect 5776 14028 7932 14056
rect 5776 14016 5782 14028
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 9398 14016 9404 14068
rect 9456 14056 9462 14068
rect 9677 14059 9735 14065
rect 9677 14056 9689 14059
rect 9456 14028 9689 14056
rect 9456 14016 9462 14028
rect 9677 14025 9689 14028
rect 9723 14025 9735 14059
rect 9677 14019 9735 14025
rect 9766 14016 9772 14068
rect 9824 14016 9830 14068
rect 11149 14059 11207 14065
rect 10520 14028 11100 14056
rect 4982 13948 4988 14000
rect 5040 13948 5046 14000
rect 9784 13988 9812 14016
rect 9416 13960 9812 13988
rect 2682 13880 2688 13932
rect 2740 13880 2746 13932
rect 4614 13920 4620 13932
rect 2884 13892 4620 13920
rect 2884 13861 2912 13892
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 5000 13920 5028 13948
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 5000 13892 5089 13920
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5534 13880 5540 13932
rect 5592 13880 5598 13932
rect 9416 13929 9444 13960
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13920 9643 13923
rect 10520 13920 10548 14028
rect 11072 13988 11100 14028
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 11422 14056 11428 14068
rect 11195 14028 11428 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 15562 14056 15568 14068
rect 12032 14028 15568 14056
rect 12032 14016 12038 14028
rect 11514 13988 11520 14000
rect 11072 13960 11520 13988
rect 11514 13948 11520 13960
rect 11572 13948 11578 14000
rect 9631 13892 10548 13920
rect 10597 13923 10655 13929
rect 9631 13889 9643 13892
rect 9585 13883 9643 13889
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 10686 13920 10692 13932
rect 10643 13892 10692 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 13740 13929 13768 14028
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 14458 13948 14464 14000
rect 14516 13948 14522 14000
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13821 2927 13855
rect 2869 13815 2927 13821
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 3007 13824 3341 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 3329 13815 3387 13821
rect 3878 13812 3884 13864
rect 3936 13812 3942 13864
rect 9030 13812 9036 13864
rect 9088 13812 9094 13864
rect 9122 13812 9128 13864
rect 9180 13812 9186 13864
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 11054 13852 11060 13864
rect 10367 13824 11060 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 13078 13812 13084 13864
rect 13136 13812 13142 13864
rect 13633 13855 13691 13861
rect 13633 13821 13645 13855
rect 13679 13852 13691 13855
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13679 13824 14013 13852
rect 13679 13821 13691 13824
rect 13633 13815 13691 13821
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 15010 13812 15016 13864
rect 15068 13852 15074 13864
rect 15473 13855 15531 13861
rect 15473 13852 15485 13855
rect 15068 13824 15485 13852
rect 15068 13812 15074 13824
rect 2498 13676 2504 13728
rect 2556 13676 2562 13728
rect 14550 13676 14556 13728
rect 14608 13716 14614 13728
rect 15120 13716 15148 13824
rect 15473 13821 15485 13824
rect 15519 13821 15531 13855
rect 15473 13815 15531 13821
rect 14608 13688 15148 13716
rect 14608 13676 14614 13688
rect 1104 13626 16008 13648
rect 1104 13574 2813 13626
rect 2865 13574 2877 13626
rect 2929 13574 2941 13626
rect 2993 13574 3005 13626
rect 3057 13574 3069 13626
rect 3121 13574 6539 13626
rect 6591 13574 6603 13626
rect 6655 13574 6667 13626
rect 6719 13574 6731 13626
rect 6783 13574 6795 13626
rect 6847 13574 10265 13626
rect 10317 13574 10329 13626
rect 10381 13574 10393 13626
rect 10445 13574 10457 13626
rect 10509 13574 10521 13626
rect 10573 13574 13991 13626
rect 14043 13574 14055 13626
rect 14107 13574 14119 13626
rect 14171 13574 14183 13626
rect 14235 13574 14247 13626
rect 14299 13574 16008 13626
rect 1104 13552 16008 13574
rect 11054 13472 11060 13524
rect 11112 13472 11118 13524
rect 13078 13472 13084 13524
rect 13136 13512 13142 13524
rect 13357 13515 13415 13521
rect 13357 13512 13369 13515
rect 13136 13484 13369 13512
rect 13136 13472 13142 13484
rect 13357 13481 13369 13484
rect 13403 13481 13415 13515
rect 13357 13475 13415 13481
rect 11330 13404 11336 13456
rect 11388 13404 11394 13456
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13376 2099 13379
rect 2498 13376 2504 13388
rect 2087 13348 2504 13376
rect 2087 13345 2099 13348
rect 2041 13339 2099 13345
rect 2498 13336 2504 13348
rect 2556 13336 2562 13388
rect 8757 13379 8815 13385
rect 8757 13345 8769 13379
rect 8803 13376 8815 13379
rect 9674 13376 9680 13388
rect 8803 13348 9680 13376
rect 8803 13345 8815 13348
rect 8757 13339 8815 13345
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 10686 13376 10692 13388
rect 10367 13348 10692 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 10873 13379 10931 13385
rect 10873 13376 10885 13379
rect 10827 13348 10885 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 10873 13345 10885 13348
rect 10919 13345 10931 13379
rect 10873 13339 10931 13345
rect 1765 13311 1823 13317
rect 1765 13277 1777 13311
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 1780 13240 1808 13271
rect 3142 13268 3148 13320
rect 3200 13268 3206 13320
rect 3326 13268 3332 13320
rect 3384 13308 3390 13320
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 3384 13280 3801 13308
rect 3384 13268 3390 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 4338 13268 4344 13320
rect 4396 13268 4402 13320
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6972 13280 7021 13308
rect 6972 13268 6978 13280
rect 7009 13277 7021 13280
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 9766 13268 9772 13320
rect 9824 13268 9830 13320
rect 10413 13311 10471 13317
rect 10413 13277 10425 13311
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 7285 13243 7343 13249
rect 1780 13212 1992 13240
rect 1964 13184 1992 13212
rect 7285 13209 7297 13243
rect 7331 13240 7343 13243
rect 7558 13240 7564 13252
rect 7331 13212 7564 13240
rect 7331 13209 7343 13212
rect 7285 13203 7343 13209
rect 7558 13200 7564 13212
rect 7616 13200 7622 13252
rect 8294 13200 8300 13252
rect 8352 13200 8358 13252
rect 10428 13240 10456 13271
rect 10502 13268 10508 13320
rect 10560 13268 10566 13320
rect 11348 13317 11376 13404
rect 13173 13379 13231 13385
rect 13173 13345 13185 13379
rect 13219 13376 13231 13379
rect 14093 13379 14151 13385
rect 14093 13376 14105 13379
rect 13219 13348 14105 13376
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 14093 13345 14105 13348
rect 14139 13345 14151 13379
rect 14461 13379 14519 13385
rect 14461 13376 14473 13379
rect 14093 13339 14151 13345
rect 14200 13348 14473 13376
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13308 10655 13311
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 10643 13280 11345 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 14200 13308 14228 13348
rect 14461 13345 14473 13348
rect 14507 13345 14519 13379
rect 14461 13339 14519 13345
rect 14550 13336 14556 13388
rect 14608 13336 14614 13388
rect 13688 13280 14228 13308
rect 14277 13311 14335 13317
rect 13688 13268 13694 13280
rect 14277 13277 14289 13311
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13308 14427 13311
rect 14415 13280 14596 13308
rect 14415 13277 14427 13280
rect 14369 13271 14427 13277
rect 11241 13243 11299 13249
rect 10428 13212 10640 13240
rect 10612 13184 10640 13212
rect 11241 13209 11253 13243
rect 11287 13240 11299 13243
rect 11422 13240 11428 13252
rect 11287 13212 11428 13240
rect 11287 13209 11299 13212
rect 11241 13203 11299 13209
rect 11422 13200 11428 13212
rect 11480 13200 11486 13252
rect 13541 13243 13599 13249
rect 13541 13209 13553 13243
rect 13587 13240 13599 13243
rect 13906 13240 13912 13252
rect 13587 13212 13912 13240
rect 13587 13209 13599 13212
rect 13541 13203 13599 13209
rect 13906 13200 13912 13212
rect 13964 13200 13970 13252
rect 1946 13132 1952 13184
rect 2004 13132 2010 13184
rect 3050 13132 3056 13184
rect 3108 13172 3114 13184
rect 3513 13175 3571 13181
rect 3513 13172 3525 13175
rect 3108 13144 3525 13172
rect 3108 13132 3114 13144
rect 3513 13141 3525 13144
rect 3559 13172 3571 13175
rect 3878 13172 3884 13184
rect 3559 13144 3884 13172
rect 3559 13141 3571 13144
rect 3513 13135 3571 13141
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 9214 13132 9220 13184
rect 9272 13132 9278 13184
rect 10594 13132 10600 13184
rect 10652 13132 10658 13184
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 14292 13172 14320 13271
rect 14568 13184 14596 13280
rect 13780 13144 14320 13172
rect 13780 13132 13786 13144
rect 14550 13132 14556 13184
rect 14608 13132 14614 13184
rect 1104 13082 16008 13104
rect 1104 13030 3473 13082
rect 3525 13030 3537 13082
rect 3589 13030 3601 13082
rect 3653 13030 3665 13082
rect 3717 13030 3729 13082
rect 3781 13030 7199 13082
rect 7251 13030 7263 13082
rect 7315 13030 7327 13082
rect 7379 13030 7391 13082
rect 7443 13030 7455 13082
rect 7507 13030 10925 13082
rect 10977 13030 10989 13082
rect 11041 13030 11053 13082
rect 11105 13030 11117 13082
rect 11169 13030 11181 13082
rect 11233 13030 14651 13082
rect 14703 13030 14715 13082
rect 14767 13030 14779 13082
rect 14831 13030 14843 13082
rect 14895 13030 14907 13082
rect 14959 13030 16008 13082
rect 1104 13008 16008 13030
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 3418 12968 3424 12980
rect 3200 12940 3424 12968
rect 3200 12928 3206 12940
rect 3418 12928 3424 12940
rect 3476 12928 3482 12980
rect 3605 12971 3663 12977
rect 3605 12937 3617 12971
rect 3651 12968 3663 12971
rect 3651 12940 4384 12968
rect 3651 12937 3663 12940
rect 3605 12931 3663 12937
rect 2866 12860 2872 12912
rect 2924 12860 2930 12912
rect 4356 12844 4384 12940
rect 4982 12928 4988 12980
rect 5040 12968 5046 12980
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 5040 12940 5181 12968
rect 5040 12928 5046 12940
rect 5169 12937 5181 12940
rect 5215 12937 5227 12971
rect 5169 12931 5227 12937
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 7745 12971 7803 12977
rect 7745 12968 7757 12971
rect 7616 12940 7757 12968
rect 7616 12928 7622 12940
rect 7745 12937 7757 12940
rect 7791 12937 7803 12971
rect 7745 12931 7803 12937
rect 9030 12928 9036 12980
rect 9088 12928 9094 12980
rect 9214 12968 9220 12980
rect 9140 12940 9220 12968
rect 5261 12903 5319 12909
rect 5261 12900 5273 12903
rect 5092 12872 5273 12900
rect 5092 12844 5120 12872
rect 5261 12869 5273 12872
rect 5307 12900 5319 12903
rect 8297 12903 8355 12909
rect 8297 12900 8309 12903
rect 5307 12872 6040 12900
rect 5307 12869 5319 12872
rect 5261 12863 5319 12869
rect 4338 12792 4344 12844
rect 4396 12792 4402 12844
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 1857 12767 1915 12773
rect 1857 12733 1869 12767
rect 1903 12764 1915 12767
rect 1903 12736 1992 12764
rect 1903 12733 1915 12736
rect 1857 12727 1915 12733
rect 1964 12640 1992 12736
rect 2130 12724 2136 12776
rect 2188 12724 2194 12776
rect 2682 12724 2688 12776
rect 2740 12764 2746 12776
rect 4157 12767 4215 12773
rect 4157 12764 4169 12767
rect 2740 12756 3188 12764
rect 3344 12756 4169 12764
rect 2740 12736 4169 12756
rect 2740 12724 2746 12736
rect 3160 12728 3372 12736
rect 4157 12733 4169 12736
rect 4203 12733 4215 12767
rect 4157 12727 4215 12733
rect 3878 12656 3884 12708
rect 3936 12696 3942 12708
rect 4632 12696 4660 12795
rect 4798 12792 4804 12844
rect 4856 12792 4862 12844
rect 5074 12792 5080 12844
rect 5132 12792 5138 12844
rect 5166 12792 5172 12844
rect 5224 12792 5230 12844
rect 5442 12792 5448 12844
rect 5500 12792 5506 12844
rect 6012 12841 6040 12872
rect 7944 12872 8309 12900
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12801 5779 12835
rect 5721 12795 5779 12801
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6181 12835 6239 12841
rect 6181 12801 6193 12835
rect 6227 12832 6239 12835
rect 7098 12832 7104 12844
rect 6227 12804 7104 12832
rect 6227 12801 6239 12804
rect 6181 12795 6239 12801
rect 5736 12764 5764 12795
rect 7098 12792 7104 12804
rect 7156 12792 7162 12844
rect 7944 12841 7972 12872
rect 8297 12869 8309 12872
rect 8343 12869 8355 12903
rect 9048 12900 9076 12928
rect 9140 12909 9168 12940
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 8297 12863 8355 12869
rect 8588 12872 9076 12900
rect 9125 12903 9183 12909
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8588 12841 8616 12872
rect 9125 12869 9137 12903
rect 9171 12869 9183 12903
rect 9125 12863 9183 12869
rect 10134 12860 10140 12912
rect 10192 12860 10198 12912
rect 10594 12860 10600 12912
rect 10652 12900 10658 12912
rect 13633 12903 13691 12909
rect 10652 12872 11100 12900
rect 10652 12860 10658 12872
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 8444 12804 8585 12832
rect 8444 12792 8450 12804
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 11072 12841 11100 12872
rect 13633 12869 13645 12903
rect 13679 12900 13691 12903
rect 13679 12872 13952 12900
rect 13679 12869 13691 12872
rect 13633 12863 13691 12869
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 10560 12804 10977 12832
rect 10560 12792 10566 12804
rect 5902 12764 5908 12776
rect 5736 12736 5908 12764
rect 5902 12724 5908 12736
rect 5960 12764 5966 12776
rect 6454 12764 6460 12776
rect 5960 12736 6460 12764
rect 5960 12724 5966 12736
rect 6454 12724 6460 12736
rect 6512 12764 6518 12776
rect 8113 12767 8171 12773
rect 8113 12764 8125 12767
rect 6512 12736 8125 12764
rect 6512 12724 6518 12736
rect 8113 12733 8125 12736
rect 8159 12733 8171 12767
rect 8113 12727 8171 12733
rect 8205 12767 8263 12773
rect 8205 12733 8217 12767
rect 8251 12764 8263 12767
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 8251 12736 8309 12764
rect 8251 12733 8263 12736
rect 8205 12727 8263 12733
rect 8297 12733 8309 12736
rect 8343 12764 8355 12767
rect 8343 12736 8800 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 5994 12696 6000 12708
rect 3936 12668 4660 12696
rect 5460 12668 6000 12696
rect 3936 12656 3942 12668
rect 1946 12588 1952 12640
rect 2004 12588 2010 12640
rect 2866 12588 2872 12640
rect 2924 12628 2930 12640
rect 3142 12628 3148 12640
rect 2924 12600 3148 12628
rect 2924 12588 2930 12600
rect 3142 12588 3148 12600
rect 3200 12628 3206 12640
rect 5460 12628 5488 12668
rect 5994 12656 6000 12668
rect 6052 12656 6058 12708
rect 3200 12600 5488 12628
rect 3200 12588 3206 12600
rect 5534 12588 5540 12640
rect 5592 12588 5598 12640
rect 8478 12588 8484 12640
rect 8536 12588 8542 12640
rect 8772 12628 8800 12736
rect 8846 12724 8852 12776
rect 8904 12724 8910 12776
rect 9858 12628 9864 12640
rect 8772 12600 9864 12628
rect 9858 12588 9864 12600
rect 9916 12588 9922 12640
rect 10134 12588 10140 12640
rect 10192 12628 10198 12640
rect 10594 12628 10600 12640
rect 10192 12600 10600 12628
rect 10192 12588 10198 12600
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10686 12588 10692 12640
rect 10744 12588 10750 12640
rect 10796 12628 10824 12804
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 13265 12835 13323 12841
rect 13265 12832 13277 12835
rect 13044 12804 13277 12832
rect 13044 12792 13050 12804
rect 13265 12801 13277 12804
rect 13311 12801 13323 12835
rect 13265 12795 13323 12801
rect 13446 12792 13452 12844
rect 13504 12832 13510 12844
rect 13924 12841 13952 12872
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13504 12804 13737 12832
rect 13504 12792 13510 12804
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 13725 12795 13783 12801
rect 13909 12835 13967 12841
rect 13909 12801 13921 12835
rect 13955 12832 13967 12835
rect 14550 12832 14556 12844
rect 13955 12804 14556 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 10873 12767 10931 12773
rect 10873 12733 10885 12767
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 10888 12696 10916 12727
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11204 12736 12204 12764
rect 11204 12724 11210 12736
rect 11330 12696 11336 12708
rect 10888 12668 11336 12696
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 12176 12640 12204 12736
rect 12802 12724 12808 12776
rect 12860 12724 12866 12776
rect 13170 12724 13176 12776
rect 13228 12724 13234 12776
rect 10870 12628 10876 12640
rect 10796 12600 10876 12628
rect 10870 12588 10876 12600
rect 10928 12628 10934 12640
rect 11606 12628 11612 12640
rect 10928 12600 11612 12628
rect 10928 12588 10934 12600
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 12158 12588 12164 12640
rect 12216 12588 12222 12640
rect 13354 12588 13360 12640
rect 13412 12628 13418 12640
rect 13541 12631 13599 12637
rect 13541 12628 13553 12631
rect 13412 12600 13553 12628
rect 13412 12588 13418 12600
rect 13541 12597 13553 12600
rect 13587 12597 13599 12631
rect 13541 12591 13599 12597
rect 13814 12588 13820 12640
rect 13872 12588 13878 12640
rect 1104 12538 16008 12560
rect 1104 12486 2813 12538
rect 2865 12486 2877 12538
rect 2929 12486 2941 12538
rect 2993 12486 3005 12538
rect 3057 12486 3069 12538
rect 3121 12486 6539 12538
rect 6591 12486 6603 12538
rect 6655 12486 6667 12538
rect 6719 12486 6731 12538
rect 6783 12486 6795 12538
rect 6847 12486 10265 12538
rect 10317 12486 10329 12538
rect 10381 12486 10393 12538
rect 10445 12486 10457 12538
rect 10509 12486 10521 12538
rect 10573 12486 13991 12538
rect 14043 12486 14055 12538
rect 14107 12486 14119 12538
rect 14171 12486 14183 12538
rect 14235 12486 14247 12538
rect 14299 12486 16008 12538
rect 1104 12464 16008 12486
rect 6546 12384 6552 12436
rect 6604 12384 6610 12436
rect 9769 12427 9827 12433
rect 9769 12393 9781 12427
rect 9815 12424 9827 12427
rect 9858 12424 9864 12436
rect 9815 12396 9864 12424
rect 9815 12393 9827 12396
rect 9769 12387 9827 12393
rect 9858 12384 9864 12396
rect 9916 12424 9922 12436
rect 9953 12427 10011 12433
rect 9953 12424 9965 12427
rect 9916 12396 9965 12424
rect 9916 12384 9922 12396
rect 9953 12393 9965 12396
rect 9999 12393 10011 12427
rect 11698 12424 11704 12436
rect 9953 12387 10011 12393
rect 11256 12396 11704 12424
rect 6641 12359 6699 12365
rect 6641 12325 6653 12359
rect 6687 12356 6699 12359
rect 7006 12356 7012 12368
rect 6687 12328 7012 12356
rect 6687 12325 6699 12328
rect 6641 12319 6699 12325
rect 7006 12316 7012 12328
rect 7064 12316 7070 12368
rect 9217 12359 9275 12365
rect 9217 12325 9229 12359
rect 9263 12356 9275 12359
rect 9263 12328 9812 12356
rect 9263 12325 9275 12328
rect 9217 12319 9275 12325
rect 9784 12300 9812 12328
rect 3605 12291 3663 12297
rect 3605 12257 3617 12291
rect 3651 12288 3663 12291
rect 3878 12288 3884 12300
rect 3651 12260 3884 12288
rect 3651 12257 3663 12260
rect 3605 12251 3663 12257
rect 3878 12248 3884 12260
rect 3936 12288 3942 12300
rect 3973 12291 4031 12297
rect 3973 12288 3985 12291
rect 3936 12260 3985 12288
rect 3936 12248 3942 12260
rect 3973 12257 3985 12260
rect 4019 12257 4031 12291
rect 8021 12291 8079 12297
rect 8021 12288 8033 12291
rect 3973 12251 4031 12257
rect 6564 12260 8033 12288
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12189 1915 12223
rect 1857 12183 1915 12189
rect 1872 12152 1900 12183
rect 5166 12180 5172 12232
rect 5224 12180 5230 12232
rect 5258 12180 5264 12232
rect 5316 12180 5322 12232
rect 6178 12180 6184 12232
rect 6236 12180 6242 12232
rect 6564 12229 6592 12260
rect 8021 12257 8033 12260
rect 8067 12288 8079 12291
rect 8110 12288 8116 12300
rect 8067 12260 8116 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 9766 12248 9772 12300
rect 9824 12248 9830 12300
rect 9861 12291 9919 12297
rect 9861 12257 9873 12291
rect 9907 12288 9919 12291
rect 10134 12288 10140 12300
rect 9907 12260 10140 12288
rect 9907 12257 9919 12260
rect 9861 12251 9919 12257
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10505 12291 10563 12297
rect 10505 12257 10517 12291
rect 10551 12257 10563 12291
rect 10505 12251 10563 12257
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 2133 12155 2191 12161
rect 1872 12124 1992 12152
rect 1964 12096 1992 12124
rect 2133 12121 2145 12155
rect 2179 12121 2191 12155
rect 3418 12152 3424 12164
rect 3358 12124 3424 12152
rect 2133 12115 2191 12121
rect 1946 12044 1952 12096
rect 2004 12044 2010 12096
rect 2148 12084 2176 12115
rect 3418 12112 3424 12124
rect 3476 12152 3482 12164
rect 3970 12152 3976 12164
rect 3476 12124 3976 12152
rect 3476 12112 3482 12124
rect 3970 12112 3976 12124
rect 4028 12112 4034 12164
rect 5184 12152 5212 12180
rect 6564 12152 6592 12183
rect 7558 12180 7564 12232
rect 7616 12180 7622 12232
rect 7650 12180 7656 12232
rect 7708 12180 7714 12232
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 5184 12124 6592 12152
rect 6825 12155 6883 12161
rect 6825 12121 6837 12155
rect 6871 12152 6883 12155
rect 7742 12152 7748 12164
rect 6871 12124 7748 12152
rect 6871 12121 6883 12124
rect 6825 12115 6883 12121
rect 7742 12112 7748 12124
rect 7800 12112 7806 12164
rect 7929 12155 7987 12161
rect 7929 12121 7941 12155
rect 7975 12121 7987 12155
rect 8312 12152 8340 12183
rect 8478 12180 8484 12232
rect 8536 12180 8542 12232
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9342 12223 9400 12229
rect 9342 12220 9354 12223
rect 9180 12192 9354 12220
rect 9180 12180 9186 12192
rect 9342 12189 9354 12192
rect 9388 12220 9400 12223
rect 9388 12192 9628 12220
rect 9388 12189 9400 12192
rect 9342 12183 9400 12189
rect 9600 12152 9628 12192
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10520 12220 10548 12251
rect 10778 12248 10784 12300
rect 10836 12248 10842 12300
rect 10870 12220 10876 12232
rect 9732 12192 10548 12220
rect 10704 12192 10876 12220
rect 9732 12180 9738 12192
rect 10594 12152 10600 12164
rect 8312 12124 8616 12152
rect 9600 12124 10600 12152
rect 7929 12115 7987 12121
rect 4522 12084 4528 12096
rect 2148 12056 4528 12084
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 4614 12044 4620 12096
rect 4672 12044 4678 12096
rect 4706 12044 4712 12096
rect 4764 12044 4770 12096
rect 5074 12044 5080 12096
rect 5132 12084 5138 12096
rect 5537 12087 5595 12093
rect 5537 12084 5549 12087
rect 5132 12056 5549 12084
rect 5132 12044 5138 12056
rect 5537 12053 5549 12056
rect 5583 12053 5595 12087
rect 5537 12047 5595 12053
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6788 12056 6929 12084
rect 6788 12044 6794 12056
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 7944 12084 7972 12115
rect 8588 12096 8616 12124
rect 10594 12112 10600 12124
rect 10652 12112 10658 12164
rect 8202 12084 8208 12096
rect 7944 12056 8208 12084
rect 6917 12047 6975 12053
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 9401 12087 9459 12093
rect 9401 12084 9413 12087
rect 8628 12056 9413 12084
rect 8628 12044 8634 12056
rect 9401 12053 9413 12056
rect 9447 12084 9459 12087
rect 10704 12084 10732 12192
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 11146 12180 11152 12232
rect 11204 12180 11210 12232
rect 11256 12229 11284 12396
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 12158 12384 12164 12436
rect 12216 12424 12222 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 12216 12396 13645 12424
rect 12216 12384 12222 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 12802 12316 12808 12368
rect 12860 12356 12866 12368
rect 13081 12359 13139 12365
rect 13081 12356 13093 12359
rect 12860 12328 13093 12356
rect 12860 12316 12866 12328
rect 13081 12325 13093 12328
rect 13127 12325 13139 12359
rect 13081 12319 13139 12325
rect 11974 12288 11980 12300
rect 11348 12260 11980 12288
rect 11348 12229 11376 12260
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11333 12223 11391 12229
rect 11333 12189 11345 12223
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 11348 12152 11376 12183
rect 12710 12180 12716 12232
rect 12768 12180 12774 12232
rect 13354 12180 13360 12232
rect 13412 12180 13418 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 13538 12220 13544 12232
rect 13495 12192 13544 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 14185 12223 14243 12229
rect 14185 12220 14197 12223
rect 13771 12192 14197 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 14185 12189 14197 12192
rect 14231 12189 14243 12223
rect 14185 12183 14243 12189
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 14737 12223 14795 12229
rect 14737 12220 14749 12223
rect 14608 12192 14749 12220
rect 14608 12180 14614 12192
rect 14737 12189 14749 12192
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 10796 12124 11376 12152
rect 11609 12155 11667 12161
rect 10796 12096 10824 12124
rect 11609 12121 11621 12155
rect 11655 12121 11667 12155
rect 11609 12115 11667 12121
rect 9447 12056 10732 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 10778 12044 10784 12096
rect 10836 12044 10842 12096
rect 11057 12087 11115 12093
rect 11057 12053 11069 12087
rect 11103 12084 11115 12087
rect 11624 12084 11652 12115
rect 11698 12112 11704 12164
rect 11756 12112 11762 12164
rect 13096 12124 13860 12152
rect 11103 12056 11652 12084
rect 11716 12084 11744 12112
rect 13096 12084 13124 12124
rect 13832 12096 13860 12124
rect 11716 12056 13124 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 13170 12044 13176 12096
rect 13228 12044 13234 12096
rect 13814 12044 13820 12096
rect 13872 12044 13878 12096
rect 1104 11994 16008 12016
rect 1104 11942 3473 11994
rect 3525 11942 3537 11994
rect 3589 11942 3601 11994
rect 3653 11942 3665 11994
rect 3717 11942 3729 11994
rect 3781 11942 7199 11994
rect 7251 11942 7263 11994
rect 7315 11942 7327 11994
rect 7379 11942 7391 11994
rect 7443 11942 7455 11994
rect 7507 11942 10925 11994
rect 10977 11942 10989 11994
rect 11041 11942 11053 11994
rect 11105 11942 11117 11994
rect 11169 11942 11181 11994
rect 11233 11942 14651 11994
rect 14703 11942 14715 11994
rect 14767 11942 14779 11994
rect 14831 11942 14843 11994
rect 14895 11942 14907 11994
rect 14959 11942 16008 11994
rect 1104 11920 16008 11942
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 2188 11852 2421 11880
rect 2188 11840 2194 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 3878 11840 3884 11892
rect 3936 11840 3942 11892
rect 6178 11840 6184 11892
rect 6236 11840 6242 11892
rect 7742 11840 7748 11892
rect 7800 11880 7806 11892
rect 7800 11852 8064 11880
rect 7800 11840 7806 11852
rect 3234 11772 3240 11824
rect 3292 11812 3298 11824
rect 3510 11812 3516 11824
rect 3292 11784 3516 11812
rect 3292 11772 3298 11784
rect 3510 11772 3516 11784
rect 3568 11772 3574 11824
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11744 2651 11747
rect 2682 11744 2688 11756
rect 2639 11716 2688 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 3326 11744 3332 11756
rect 2915 11716 3332 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 3896 11744 3924 11840
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 6822 11812 6828 11824
rect 4028 11784 5198 11812
rect 6472 11784 6828 11812
rect 4028 11772 4034 11784
rect 4430 11744 4436 11756
rect 3835 11716 3924 11744
rect 3988 11716 4436 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 3234 11636 3240 11688
rect 3292 11636 3298 11688
rect 3988 11676 4016 11716
rect 4430 11704 4436 11716
rect 4488 11704 4494 11756
rect 3436 11648 4016 11676
rect 4065 11679 4123 11685
rect 1946 11568 1952 11620
rect 2004 11608 2010 11620
rect 3436 11608 3464 11648
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 4246 11676 4252 11688
rect 4111 11648 4252 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 4338 11636 4344 11688
rect 4396 11636 4402 11688
rect 4706 11636 4712 11688
rect 4764 11636 4770 11688
rect 5442 11636 5448 11688
rect 5500 11676 5506 11688
rect 6472 11685 6500 11784
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 8036 11744 8064 11852
rect 8202 11840 8208 11892
rect 8260 11840 8266 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 10045 11883 10103 11889
rect 10045 11880 10057 11883
rect 8536 11852 10057 11880
rect 8536 11840 8542 11852
rect 10045 11849 10057 11852
rect 10091 11849 10103 11883
rect 10045 11843 10103 11849
rect 10134 11840 10140 11892
rect 10192 11840 10198 11892
rect 13170 11840 13176 11892
rect 13228 11840 13234 11892
rect 8220 11812 8248 11840
rect 8297 11815 8355 11821
rect 8297 11812 8309 11815
rect 8220 11784 8309 11812
rect 8297 11781 8309 11784
rect 8343 11781 8355 11815
rect 8297 11775 8355 11781
rect 10152 11753 10180 11840
rect 13081 11815 13139 11821
rect 13081 11781 13093 11815
rect 13127 11812 13139 11815
rect 13188 11812 13216 11840
rect 13127 11784 13216 11812
rect 13127 11781 13139 11784
rect 13081 11775 13139 11781
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 7866 11716 7972 11744
rect 8036 11716 8493 11744
rect 6457 11679 6515 11685
rect 6457 11676 6469 11679
rect 5500 11648 6469 11676
rect 5500 11636 5506 11648
rect 6457 11645 6469 11648
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 6730 11636 6736 11688
rect 6788 11636 6794 11688
rect 2004 11580 3464 11608
rect 2004 11568 2010 11580
rect 3510 11568 3516 11620
rect 3568 11568 3574 11620
rect 3697 11611 3755 11617
rect 3697 11577 3709 11611
rect 3743 11608 3755 11611
rect 3786 11608 3792 11620
rect 3743 11580 3792 11608
rect 3743 11577 3755 11580
rect 3697 11571 3755 11577
rect 3786 11568 3792 11580
rect 3844 11568 3850 11620
rect 4356 11608 4384 11636
rect 4172 11580 4384 11608
rect 7944 11608 7972 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 10137 11747 10195 11753
rect 10137 11713 10149 11747
rect 10183 11713 10195 11747
rect 10137 11707 10195 11713
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 8018 11636 8024 11688
rect 8076 11676 8082 11688
rect 8680 11676 8708 11707
rect 8076 11648 8708 11676
rect 11517 11679 11575 11685
rect 8076 11636 8082 11648
rect 11517 11645 11529 11679
rect 11563 11676 11575 11679
rect 11698 11676 11704 11688
rect 11563 11648 11704 11676
rect 11563 11645 11575 11648
rect 11517 11639 11575 11645
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 7944 11580 8524 11608
rect 2777 11543 2835 11549
rect 2777 11509 2789 11543
rect 2823 11540 2835 11543
rect 3142 11540 3148 11552
rect 2823 11512 3148 11540
rect 2823 11509 2835 11512
rect 2777 11503 2835 11509
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 3528 11540 3556 11568
rect 3878 11540 3884 11552
rect 3528 11512 3884 11540
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4172 11549 4200 11580
rect 8496 11552 8524 11580
rect 8570 11568 8576 11620
rect 8628 11568 8634 11620
rect 11606 11568 11612 11620
rect 11664 11568 11670 11620
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 4120 11512 4169 11540
rect 4120 11500 4126 11512
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 4338 11500 4344 11552
rect 4396 11500 4402 11552
rect 8478 11500 8484 11552
rect 8536 11500 8542 11552
rect 11900 11540 11928 11707
rect 11974 11704 11980 11756
rect 12032 11744 12038 11756
rect 12802 11744 12808 11756
rect 12032 11716 12808 11744
rect 12032 11704 12038 11716
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 14366 11744 14372 11756
rect 14214 11716 14372 11744
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11676 12127 11679
rect 14550 11676 14556 11688
rect 12115 11648 14556 11676
rect 12115 11645 12127 11648
rect 12069 11639 12127 11645
rect 14550 11636 14556 11648
rect 14608 11636 14614 11688
rect 13538 11540 13544 11552
rect 11900 11512 13544 11540
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 1104 11450 16008 11472
rect 1104 11398 2813 11450
rect 2865 11398 2877 11450
rect 2929 11398 2941 11450
rect 2993 11398 3005 11450
rect 3057 11398 3069 11450
rect 3121 11398 6539 11450
rect 6591 11398 6603 11450
rect 6655 11398 6667 11450
rect 6719 11398 6731 11450
rect 6783 11398 6795 11450
rect 6847 11398 10265 11450
rect 10317 11398 10329 11450
rect 10381 11398 10393 11450
rect 10445 11398 10457 11450
rect 10509 11398 10521 11450
rect 10573 11398 13991 11450
rect 14043 11398 14055 11450
rect 14107 11398 14119 11450
rect 14171 11398 14183 11450
rect 14235 11398 14247 11450
rect 14299 11398 16008 11450
rect 1104 11376 16008 11398
rect 3326 11296 3332 11348
rect 3384 11336 3390 11348
rect 3881 11339 3939 11345
rect 3384 11308 3740 11336
rect 3384 11296 3390 11308
rect 3234 11228 3240 11280
rect 3292 11268 3298 11280
rect 3712 11268 3740 11308
rect 3881 11305 3893 11339
rect 3927 11336 3939 11339
rect 4154 11336 4160 11348
rect 3927 11308 4160 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4246 11296 4252 11348
rect 4304 11296 4310 11348
rect 4338 11296 4344 11348
rect 4396 11296 4402 11348
rect 4430 11296 4436 11348
rect 4488 11296 4494 11348
rect 4522 11296 4528 11348
rect 4580 11296 4586 11348
rect 4893 11339 4951 11345
rect 4893 11305 4905 11339
rect 4939 11336 4951 11339
rect 5258 11336 5264 11348
rect 4939 11308 5264 11336
rect 4939 11305 4951 11308
rect 4893 11299 4951 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 5432 11339 5490 11345
rect 5432 11305 5444 11339
rect 5478 11336 5490 11339
rect 5534 11336 5540 11348
rect 5478 11308 5540 11336
rect 5478 11305 5490 11308
rect 5432 11299 5490 11305
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 7745 11339 7803 11345
rect 7745 11336 7757 11339
rect 7616 11308 7757 11336
rect 7616 11296 7622 11308
rect 7745 11305 7757 11308
rect 7791 11305 7803 11339
rect 7745 11299 7803 11305
rect 8110 11296 8116 11348
rect 8168 11296 8174 11348
rect 8202 11296 8208 11348
rect 8260 11296 8266 11348
rect 3970 11268 3976 11280
rect 3292 11240 3648 11268
rect 3712 11240 3976 11268
rect 3292 11228 3298 11240
rect 3620 11209 3648 11240
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 2961 11203 3019 11209
rect 2961 11169 2973 11203
rect 3007 11200 3019 11203
rect 3513 11203 3571 11209
rect 3007 11172 3464 11200
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 2869 11135 2927 11141
rect 2869 11132 2881 11135
rect 2792 11104 2881 11132
rect 2792 11064 2820 11104
rect 2869 11101 2881 11104
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3329 11135 3387 11141
rect 3099 11104 3280 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3252 11076 3280 11104
rect 3329 11101 3341 11135
rect 3375 11101 3387 11135
rect 3329 11095 3387 11101
rect 3145 11067 3203 11073
rect 3145 11064 3157 11067
rect 2792 11036 3157 11064
rect 2792 11008 2820 11036
rect 3145 11033 3157 11036
rect 3191 11033 3203 11067
rect 3145 11027 3203 11033
rect 3234 11024 3240 11076
rect 3292 11024 3298 11076
rect 2774 10956 2780 11008
rect 2832 10956 2838 11008
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 3344 10996 3372 11095
rect 3436 11064 3464 11172
rect 3513 11169 3525 11203
rect 3559 11169 3571 11203
rect 3513 11163 3571 11169
rect 3605 11203 3663 11209
rect 3605 11169 3617 11203
rect 3651 11200 3663 11203
rect 4062 11200 4068 11220
rect 3651 11172 4068 11200
rect 3651 11169 3663 11172
rect 3605 11163 3663 11169
rect 4062 11168 4068 11172
rect 4120 11168 4126 11220
rect 4065 11163 4123 11168
rect 3528 11132 3556 11163
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3528 11104 3801 11132
rect 3789 11101 3801 11104
rect 3835 11132 3847 11135
rect 4264 11132 4292 11296
rect 4356 11200 4384 11296
rect 4448 11268 4476 11296
rect 4448 11240 5212 11268
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4356 11172 4445 11200
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4798 11160 4804 11212
rect 4856 11160 4862 11212
rect 5184 11209 5212 11240
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 8018 11268 8024 11280
rect 7064 11240 8024 11268
rect 7064 11228 7070 11240
rect 8018 11228 8024 11240
rect 8076 11228 8082 11280
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 5534 11200 5540 11212
rect 5215 11172 5540 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5994 11160 6000 11212
rect 6052 11200 6058 11212
rect 6052 11172 6684 11200
rect 6052 11160 6058 11172
rect 3835 11104 4292 11132
rect 3835 11101 3847 11104
rect 3789 11095 3847 11101
rect 4338 11092 4344 11144
rect 4396 11092 4402 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4632 11064 4660 11095
rect 4706 11092 4712 11144
rect 4764 11092 4770 11144
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5000 11064 5028 11095
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 3436 11036 5028 11064
rect 6656 11064 6684 11172
rect 7742 11160 7748 11212
rect 7800 11160 7806 11212
rect 8128 11209 8156 11296
rect 8220 11209 8248 11296
rect 12710 11268 12716 11280
rect 11900 11240 12716 11268
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 9674 11160 9680 11212
rect 9732 11160 9738 11212
rect 9953 11203 10011 11209
rect 9953 11169 9965 11203
rect 9999 11200 10011 11203
rect 11330 11200 11336 11212
rect 9999 11172 11336 11200
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 11330 11160 11336 11172
rect 11388 11160 11394 11212
rect 11425 11203 11483 11209
rect 11425 11169 11437 11203
rect 11471 11200 11483 11203
rect 11790 11200 11796 11212
rect 11471 11172 11796 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 11790 11160 11796 11172
rect 11848 11160 11854 11212
rect 7760 11132 7788 11160
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7760 11104 7941 11132
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8444 11104 8953 11132
rect 8444 11092 8450 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9490 11092 9496 11144
rect 9548 11092 9554 11144
rect 11514 11132 11520 11144
rect 11086 11104 11520 11132
rect 11514 11092 11520 11104
rect 11572 11132 11578 11144
rect 11900 11132 11928 11240
rect 12710 11228 12716 11240
rect 12768 11268 12774 11280
rect 13446 11268 13452 11280
rect 12768 11240 13452 11268
rect 12768 11228 12774 11240
rect 13446 11228 13452 11240
rect 13504 11228 13510 11280
rect 13538 11228 13544 11280
rect 13596 11268 13602 11280
rect 13817 11271 13875 11277
rect 13817 11268 13829 11271
rect 13596 11240 13829 11268
rect 13596 11228 13602 11240
rect 13817 11237 13829 11240
rect 13863 11268 13875 11271
rect 13863 11240 14504 11268
rect 13863 11237 13875 11240
rect 13817 11231 13875 11237
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11200 12587 11203
rect 12618 11200 12624 11212
rect 12575 11172 12624 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 13722 11200 13728 11212
rect 13648 11172 13728 11200
rect 12360 11134 12480 11142
rect 12713 11135 12771 11141
rect 12360 11132 12572 11134
rect 12713 11132 12725 11135
rect 11572 11104 11928 11132
rect 12268 11114 12725 11132
rect 12268 11104 12388 11114
rect 12452 11106 12725 11114
rect 12544 11104 12725 11106
rect 11572 11092 11578 11104
rect 8478 11064 8484 11076
rect 6656 11050 8484 11064
rect 6670 11036 8484 11050
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 3016 10968 3372 10996
rect 4065 10999 4123 11005
rect 3016 10956 3022 10968
rect 4065 10965 4077 10999
rect 4111 10996 4123 10999
rect 4246 10996 4252 11008
rect 4111 10968 4252 10996
rect 4111 10965 4123 10968
rect 4065 10959 4123 10965
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 5350 10956 5356 11008
rect 5408 10996 5414 11008
rect 6917 10999 6975 11005
rect 6917 10996 6929 10999
rect 5408 10968 6929 10996
rect 5408 10956 5414 10968
rect 6917 10965 6929 10968
rect 6963 10996 6975 10999
rect 7650 10996 7656 11008
rect 6963 10968 7656 10996
rect 6963 10965 6975 10968
rect 6917 10959 6975 10965
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 11422 10996 11428 11008
rect 10652 10968 11428 10996
rect 10652 10956 10658 10968
rect 11422 10956 11428 10968
rect 11480 10996 11486 11008
rect 12268 10996 12296 11104
rect 12713 11101 12725 11104
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 12820 11064 12848 11095
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 13648 11141 13676 11172
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 14476 11209 14504 11240
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 13449 11135 13507 11141
rect 13449 11132 13461 11135
rect 13412 11104 13461 11132
rect 13412 11092 13418 11104
rect 13449 11101 13461 11104
rect 13495 11101 13507 11135
rect 13449 11095 13507 11101
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11132 13691 11135
rect 13885 11135 13943 11141
rect 13885 11132 13897 11135
rect 13679 11104 13897 11132
rect 13679 11101 13691 11104
rect 13633 11095 13691 11101
rect 13885 11101 13897 11104
rect 13931 11101 13943 11135
rect 13885 11095 13943 11101
rect 14553 11135 14611 11141
rect 14553 11101 14565 11135
rect 14599 11132 14611 11135
rect 15010 11132 15016 11144
rect 14599 11104 15016 11132
rect 14599 11101 14611 11104
rect 14553 11095 14611 11101
rect 12360 11036 12848 11064
rect 13464 11064 13492 11095
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 13722 11064 13728 11076
rect 13464 11036 13728 11064
rect 12360 11008 12388 11036
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 14093 11067 14151 11073
rect 14093 11064 14105 11067
rect 13832 11036 14105 11064
rect 11480 10968 12296 10996
rect 11480 10956 11486 10968
rect 12342 10956 12348 11008
rect 12400 10956 12406 11008
rect 12434 10956 12440 11008
rect 12492 10956 12498 11008
rect 12526 10956 12532 11008
rect 12584 10956 12590 11008
rect 13541 10999 13599 11005
rect 13541 10965 13553 10999
rect 13587 10996 13599 10999
rect 13832 10996 13860 11036
rect 14093 11033 14105 11036
rect 14139 11064 14151 11067
rect 14139 11036 14320 11064
rect 14139 11033 14151 11036
rect 14093 11027 14151 11033
rect 13587 10968 13860 10996
rect 14292 10996 14320 11036
rect 14366 11024 14372 11076
rect 14424 11064 14430 11076
rect 14829 11067 14887 11073
rect 14829 11064 14841 11067
rect 14424 11036 14841 11064
rect 14424 11024 14430 11036
rect 14829 11033 14841 11036
rect 14875 11033 14887 11067
rect 14829 11027 14887 11033
rect 15197 11067 15255 11073
rect 15197 11033 15209 11067
rect 15243 11064 15255 11067
rect 15378 11064 15384 11076
rect 15243 11036 15384 11064
rect 15243 11033 15255 11036
rect 15197 11027 15255 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 14458 10996 14464 11008
rect 14292 10968 14464 10996
rect 13587 10965 13599 10968
rect 13541 10959 13599 10965
rect 14458 10956 14464 10968
rect 14516 10956 14522 11008
rect 14550 10956 14556 11008
rect 14608 10996 14614 11008
rect 14737 10999 14795 11005
rect 14737 10996 14749 10999
rect 14608 10968 14749 10996
rect 14608 10956 14614 10968
rect 14737 10965 14749 10968
rect 14783 10965 14795 10999
rect 14737 10959 14795 10965
rect 1104 10906 16008 10928
rect 1104 10854 3473 10906
rect 3525 10854 3537 10906
rect 3589 10854 3601 10906
rect 3653 10854 3665 10906
rect 3717 10854 3729 10906
rect 3781 10854 7199 10906
rect 7251 10854 7263 10906
rect 7315 10854 7327 10906
rect 7379 10854 7391 10906
rect 7443 10854 7455 10906
rect 7507 10854 10925 10906
rect 10977 10854 10989 10906
rect 11041 10854 11053 10906
rect 11105 10854 11117 10906
rect 11169 10854 11181 10906
rect 11233 10854 14651 10906
rect 14703 10854 14715 10906
rect 14767 10854 14779 10906
rect 14831 10854 14843 10906
rect 14895 10854 14907 10906
rect 14959 10854 16008 10906
rect 1104 10832 16008 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 3142 10792 3148 10804
rect 1627 10764 3148 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 8665 10795 8723 10801
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 9490 10792 9496 10804
rect 8711 10764 9496 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10778 10792 10784 10804
rect 9732 10764 10784 10792
rect 9732 10752 9738 10764
rect 10778 10752 10784 10764
rect 10836 10792 10842 10804
rect 10873 10795 10931 10801
rect 10873 10792 10885 10795
rect 10836 10764 10885 10792
rect 10836 10752 10842 10764
rect 10873 10761 10885 10764
rect 10919 10761 10931 10795
rect 10873 10755 10931 10761
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11388 10764 11529 10792
rect 11388 10752 11394 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11664 10764 11713 10792
rect 11664 10752 11670 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 11701 10755 11759 10761
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12860 10764 14964 10792
rect 12860 10752 12866 10764
rect 2866 10684 2872 10736
rect 2924 10684 2930 10736
rect 8478 10724 8484 10736
rect 8418 10696 8484 10724
rect 8478 10684 8484 10696
rect 8536 10724 8542 10736
rect 8757 10727 8815 10733
rect 8757 10724 8769 10727
rect 8536 10696 8769 10724
rect 8536 10684 8542 10696
rect 8757 10693 8769 10696
rect 8803 10693 8815 10727
rect 14366 10724 14372 10736
rect 14214 10696 14372 10724
rect 8757 10687 8815 10693
rect 14366 10684 14372 10696
rect 14424 10684 14430 10736
rect 14550 10684 14556 10736
rect 14608 10724 14614 10736
rect 14645 10727 14703 10733
rect 14645 10724 14657 10727
rect 14608 10696 14657 10724
rect 14608 10684 14614 10696
rect 14645 10693 14657 10696
rect 14691 10693 14703 10727
rect 14645 10687 14703 10693
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 4212 10628 4721 10656
rect 4212 10616 4218 10628
rect 4709 10625 4721 10628
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 4982 10616 4988 10668
rect 5040 10616 5046 10668
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10656 5227 10659
rect 5350 10656 5356 10668
rect 5215 10628 5356 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 5592 10628 6929 10656
rect 5592 10616 5598 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 9125 10659 9183 10665
rect 9125 10625 9137 10659
rect 9171 10656 9183 10659
rect 9214 10656 9220 10668
rect 9171 10628 9220 10656
rect 9171 10625 9183 10628
rect 9125 10619 9183 10625
rect 9214 10616 9220 10628
rect 9272 10616 9278 10668
rect 9582 10616 9588 10668
rect 9640 10616 9646 10668
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 11655 10659 11713 10665
rect 11480 10646 11560 10656
rect 11655 10646 11667 10659
rect 11480 10628 11667 10646
rect 11480 10616 11486 10628
rect 11532 10625 11667 10628
rect 11701 10625 11713 10659
rect 11532 10619 11713 10625
rect 11532 10618 11685 10619
rect 11790 10616 11796 10668
rect 11848 10656 11854 10668
rect 12253 10659 12311 10665
rect 12253 10656 12265 10659
rect 11848 10628 12265 10656
rect 11848 10616 11854 10628
rect 12253 10625 12265 10628
rect 12299 10625 12311 10659
rect 12253 10619 12311 10625
rect 13630 10616 13636 10668
rect 13688 10616 13694 10668
rect 14936 10665 14964 10764
rect 15010 10752 15016 10804
rect 15068 10752 15074 10804
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10625 14979 10659
rect 14921 10619 14979 10625
rect 1946 10548 1952 10600
rect 2004 10548 2010 10600
rect 2222 10548 2228 10600
rect 2280 10548 2286 10600
rect 2958 10548 2964 10600
rect 3016 10588 3022 10600
rect 3697 10591 3755 10597
rect 3697 10588 3709 10591
rect 3016 10560 3709 10588
rect 3016 10548 3022 10560
rect 3697 10557 3709 10560
rect 3743 10588 3755 10591
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 3743 10560 4445 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 4433 10557 4445 10560
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 4448 10520 4476 10551
rect 4614 10548 4620 10600
rect 4672 10548 4678 10600
rect 7190 10548 7196 10600
rect 7248 10548 7254 10600
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12434 10588 12440 10600
rect 12207 10560 12440 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 13173 10591 13231 10597
rect 13173 10557 13185 10591
rect 13219 10588 13231 10591
rect 13648 10588 13676 10616
rect 13219 10560 13676 10588
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 15102 10548 15108 10600
rect 15160 10588 15166 10600
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 15160 10560 15577 10588
rect 15160 10548 15166 10560
rect 15565 10557 15577 10560
rect 15611 10557 15623 10591
rect 15565 10551 15623 10557
rect 12069 10523 12127 10529
rect 4448 10492 5212 10520
rect 5184 10464 5212 10492
rect 12069 10489 12081 10523
rect 12115 10520 12127 10523
rect 12618 10520 12624 10532
rect 12115 10492 12624 10520
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 3786 10412 3792 10464
rect 3844 10412 3850 10464
rect 5166 10412 5172 10464
rect 5224 10412 5230 10464
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 12342 10452 12348 10464
rect 11756 10424 12348 10452
rect 11756 10412 11762 10424
rect 12342 10412 12348 10424
rect 12400 10412 12406 10464
rect 1104 10362 16008 10384
rect 1104 10310 2813 10362
rect 2865 10310 2877 10362
rect 2929 10310 2941 10362
rect 2993 10310 3005 10362
rect 3057 10310 3069 10362
rect 3121 10310 6539 10362
rect 6591 10310 6603 10362
rect 6655 10310 6667 10362
rect 6719 10310 6731 10362
rect 6783 10310 6795 10362
rect 6847 10310 10265 10362
rect 10317 10310 10329 10362
rect 10381 10310 10393 10362
rect 10445 10310 10457 10362
rect 10509 10310 10521 10362
rect 10573 10310 13991 10362
rect 14043 10310 14055 10362
rect 14107 10310 14119 10362
rect 14171 10310 14183 10362
rect 14235 10310 14247 10362
rect 14299 10310 16008 10362
rect 1104 10288 16008 10310
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2280 10220 2789 10248
rect 2280 10208 2286 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 2777 10211 2835 10217
rect 3786 10208 3792 10260
rect 3844 10208 3850 10260
rect 5534 10208 5540 10260
rect 5592 10208 5598 10260
rect 7098 10208 7104 10260
rect 7156 10208 7162 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7248 10220 7849 10248
rect 7248 10208 7254 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 7837 10211 7895 10217
rect 12529 10251 12587 10257
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12618 10248 12624 10260
rect 12575 10220 12624 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 15010 10208 15016 10260
rect 15068 10208 15074 10260
rect 3142 10072 3148 10124
rect 3200 10112 3206 10124
rect 3421 10115 3479 10121
rect 3200 10084 3372 10112
rect 3200 10072 3206 10084
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 3344 10053 3372 10084
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 3804 10112 3832 10208
rect 13722 10140 13728 10192
rect 13780 10180 13786 10192
rect 13780 10152 14964 10180
rect 13780 10140 13786 10152
rect 3467 10084 3832 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 7650 10072 7656 10124
rect 7708 10072 7714 10124
rect 8481 10115 8539 10121
rect 8481 10112 8493 10115
rect 8036 10084 8493 10112
rect 2902 10047 2960 10053
rect 2902 10044 2914 10047
rect 2832 10016 2914 10044
rect 2832 10004 2838 10016
rect 2902 10013 2914 10016
rect 2948 10044 2960 10047
rect 3329 10047 3387 10053
rect 2948 10016 3280 10044
rect 2948 10013 2960 10016
rect 2902 10007 2960 10013
rect 3252 9976 3280 10016
rect 3329 10013 3341 10047
rect 3375 10044 3387 10047
rect 3878 10044 3884 10056
rect 3375 10016 3884 10044
rect 3375 10013 3387 10016
rect 3329 10007 3387 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 8036 10053 8064 10084
rect 8481 10081 8493 10084
rect 8527 10081 8539 10115
rect 8481 10075 8539 10081
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 9769 10115 9827 10121
rect 9769 10112 9781 10115
rect 9732 10084 9781 10112
rect 9732 10072 9738 10084
rect 9769 10081 9781 10084
rect 9815 10081 9827 10115
rect 9769 10075 9827 10081
rect 10045 10115 10103 10121
rect 10045 10081 10057 10115
rect 10091 10112 10103 10115
rect 11330 10112 11336 10124
rect 10091 10084 11336 10112
rect 10091 10081 10103 10084
rect 10045 10075 10103 10081
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11563 10084 11897 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 11885 10081 11897 10084
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 13630 10072 13636 10124
rect 13688 10072 13694 10124
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 14829 10115 14887 10121
rect 14829 10112 14841 10115
rect 13964 10084 14841 10112
rect 13964 10072 13970 10084
rect 14829 10081 14841 10084
rect 14875 10081 14887 10115
rect 14829 10075 14887 10081
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 8202 10004 8208 10056
rect 8260 10004 8266 10056
rect 8297 10047 8355 10053
rect 8297 10013 8309 10047
rect 8343 10044 8355 10047
rect 8386 10044 8392 10056
rect 8343 10016 8392 10044
rect 8343 10013 8355 10016
rect 8297 10007 8355 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 13648 10044 13676 10072
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13648 10016 14105 10044
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14936 10044 14964 10152
rect 15028 10112 15056 10208
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 15028 10084 15117 10112
rect 15105 10081 15117 10084
rect 15151 10081 15163 10115
rect 15105 10075 15163 10081
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 14936 10016 15025 10044
rect 14093 10007 14151 10013
rect 15013 10013 15025 10016
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 15197 10047 15255 10053
rect 15197 10013 15209 10047
rect 15243 10013 15255 10047
rect 15197 10007 15255 10013
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 4062 9976 4068 9988
rect 3252 9948 4068 9976
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 6914 9936 6920 9988
rect 6972 9976 6978 9988
rect 7009 9979 7067 9985
rect 7009 9976 7021 9979
rect 6972 9948 7021 9976
rect 6972 9936 6978 9948
rect 7009 9945 7021 9948
rect 7055 9976 7067 9979
rect 9582 9976 9588 9988
rect 7055 9948 9588 9976
rect 7055 9945 7067 9948
rect 7009 9939 7067 9945
rect 9582 9936 9588 9948
rect 9640 9936 9646 9988
rect 11514 9976 11520 9988
rect 11270 9948 11520 9976
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 14737 9979 14795 9985
rect 14737 9945 14749 9979
rect 14783 9976 14795 9979
rect 15212 9976 15240 10007
rect 14783 9948 15240 9976
rect 14783 9945 14795 9948
rect 14737 9939 14795 9945
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 3234 9908 3240 9920
rect 3007 9880 3240 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 3234 9868 3240 9880
rect 3292 9908 3298 9920
rect 4154 9908 4160 9920
rect 3292 9880 4160 9908
rect 3292 9868 3298 9880
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 15304 9908 15332 10007
rect 15068 9880 15332 9908
rect 15068 9868 15074 9880
rect 1104 9818 16008 9840
rect 1104 9766 3473 9818
rect 3525 9766 3537 9818
rect 3589 9766 3601 9818
rect 3653 9766 3665 9818
rect 3717 9766 3729 9818
rect 3781 9766 7199 9818
rect 7251 9766 7263 9818
rect 7315 9766 7327 9818
rect 7379 9766 7391 9818
rect 7443 9766 7455 9818
rect 7507 9766 10925 9818
rect 10977 9766 10989 9818
rect 11041 9766 11053 9818
rect 11105 9766 11117 9818
rect 11169 9766 11181 9818
rect 11233 9766 14651 9818
rect 14703 9766 14715 9818
rect 14767 9766 14779 9818
rect 14831 9766 14843 9818
rect 14895 9766 14907 9818
rect 14959 9766 16008 9818
rect 1104 9744 16008 9766
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 4249 9707 4307 9713
rect 4249 9704 4261 9707
rect 4212 9676 4261 9704
rect 4212 9664 4218 9676
rect 4249 9673 4261 9676
rect 4295 9673 4307 9707
rect 4249 9667 4307 9673
rect 11330 9664 11336 9716
rect 11388 9664 11394 9716
rect 12250 9664 12256 9716
rect 12308 9704 12314 9716
rect 12618 9704 12624 9716
rect 12308 9676 12624 9704
rect 12308 9664 12314 9676
rect 12618 9664 12624 9676
rect 12676 9664 12682 9716
rect 15102 9664 15108 9716
rect 15160 9664 15166 9716
rect 3142 9596 3148 9648
rect 3200 9636 3206 9648
rect 3513 9639 3571 9645
rect 3513 9636 3525 9639
rect 3200 9608 3525 9636
rect 3200 9596 3206 9608
rect 3513 9605 3525 9608
rect 3559 9605 3571 9639
rect 5261 9639 5319 9645
rect 5261 9636 5273 9639
rect 3513 9599 3571 9605
rect 3896 9608 5273 9636
rect 3896 9580 3924 9608
rect 5261 9605 5273 9608
rect 5307 9605 5319 9639
rect 11348 9636 11376 9664
rect 11609 9639 11667 9645
rect 11609 9636 11621 9639
rect 11348 9608 11621 9636
rect 5261 9599 5319 9605
rect 11609 9605 11621 9608
rect 11655 9605 11667 9639
rect 11609 9599 11667 9605
rect 13633 9639 13691 9645
rect 13633 9605 13645 9639
rect 13679 9636 13691 9639
rect 13906 9636 13912 9648
rect 13679 9608 13912 9636
rect 13679 9605 13691 9608
rect 13633 9599 13691 9605
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 14366 9596 14372 9648
rect 14424 9596 14430 9648
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3326 9568 3332 9580
rect 3283 9540 3332 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 3344 9432 3372 9528
rect 3804 9500 3832 9531
rect 3878 9528 3884 9580
rect 3936 9528 3942 9580
rect 3970 9528 3976 9580
rect 4028 9528 4034 9580
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4190 9571 4248 9577
rect 4190 9568 4202 9571
rect 4120 9540 4202 9568
rect 4120 9528 4126 9540
rect 4190 9537 4202 9540
rect 4236 9568 4248 9571
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4236 9540 4997 9568
rect 4236 9537 4248 9540
rect 4190 9531 4248 9537
rect 4985 9537 4997 9540
rect 5031 9537 5043 9571
rect 4985 9531 5043 9537
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 3988 9500 4016 9528
rect 3804 9472 4016 9500
rect 4614 9460 4620 9512
rect 4672 9460 4678 9512
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 4798 9500 4804 9512
rect 4755 9472 4804 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 5092 9500 5120 9531
rect 5166 9528 5172 9580
rect 5224 9528 5230 9580
rect 5442 9528 5448 9580
rect 5500 9528 5506 9580
rect 8754 9528 8760 9580
rect 8812 9528 8818 9580
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 10873 9571 10931 9577
rect 10873 9568 10885 9571
rect 10836 9540 10885 9568
rect 10836 9528 10842 9540
rect 10873 9537 10885 9540
rect 10919 9537 10931 9571
rect 10873 9531 10931 9537
rect 11241 9571 11299 9577
rect 11241 9537 11253 9571
rect 11287 9568 11299 9571
rect 11330 9568 11336 9580
rect 11287 9540 11336 9568
rect 11287 9537 11299 9540
rect 11241 9531 11299 9537
rect 11330 9528 11336 9540
rect 11388 9528 11394 9580
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9568 11851 9571
rect 11839 9540 12434 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5000 9472 5549 9500
rect 4632 9432 4660 9460
rect 5000 9432 5028 9472
rect 5537 9469 5549 9472
rect 5583 9469 5595 9503
rect 5537 9463 5595 9469
rect 9214 9460 9220 9512
rect 9272 9500 9278 9512
rect 11057 9503 11115 9509
rect 9272 9472 11008 9500
rect 9272 9460 9278 9472
rect 3344 9404 5028 9432
rect 10980 9432 11008 9472
rect 11057 9469 11069 9503
rect 11103 9500 11115 9503
rect 11698 9500 11704 9512
rect 11103 9472 11704 9500
rect 11103 9469 11115 9472
rect 11057 9463 11115 9469
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 12069 9503 12127 9509
rect 12069 9469 12081 9503
rect 12115 9500 12127 9503
rect 12250 9500 12256 9512
rect 12115 9472 12256 9500
rect 12115 9469 12127 9472
rect 12069 9463 12127 9469
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 12406 9500 12434 9540
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 12860 9540 13369 9568
rect 12860 9528 12866 9540
rect 13357 9537 13369 9540
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 12526 9500 12532 9512
rect 12406 9472 12532 9500
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 10980 9404 12434 9432
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 3786 9364 3792 9376
rect 2740 9336 3792 9364
rect 2740 9324 2746 9336
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 4062 9324 4068 9376
rect 4120 9324 4126 9376
rect 4614 9324 4620 9376
rect 4672 9324 4678 9376
rect 4890 9324 4896 9376
rect 4948 9324 4954 9376
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 10229 9367 10287 9373
rect 10229 9364 10241 9367
rect 9732 9336 10241 9364
rect 9732 9324 9738 9336
rect 10229 9333 10241 9336
rect 10275 9364 10287 9367
rect 10594 9364 10600 9376
rect 10275 9336 10600 9364
rect 10275 9333 10287 9336
rect 10229 9327 10287 9333
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 11514 9364 11520 9376
rect 11195 9336 11520 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 11514 9324 11520 9336
rect 11572 9364 11578 9376
rect 11698 9364 11704 9376
rect 11572 9336 11704 9364
rect 11572 9324 11578 9336
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 11977 9367 12035 9373
rect 11977 9364 11989 9367
rect 11940 9336 11989 9364
rect 11940 9324 11946 9336
rect 11977 9333 11989 9336
rect 12023 9333 12035 9367
rect 12406 9364 12434 9404
rect 15378 9364 15384 9376
rect 12406 9336 15384 9364
rect 11977 9327 12035 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 1104 9274 16008 9296
rect 1104 9222 2813 9274
rect 2865 9222 2877 9274
rect 2929 9222 2941 9274
rect 2993 9222 3005 9274
rect 3057 9222 3069 9274
rect 3121 9222 6539 9274
rect 6591 9222 6603 9274
rect 6655 9222 6667 9274
rect 6719 9222 6731 9274
rect 6783 9222 6795 9274
rect 6847 9222 10265 9274
rect 10317 9222 10329 9274
rect 10381 9222 10393 9274
rect 10445 9222 10457 9274
rect 10509 9222 10521 9274
rect 10573 9222 13991 9274
rect 14043 9222 14055 9274
rect 14107 9222 14119 9274
rect 14171 9222 14183 9274
rect 14235 9222 14247 9274
rect 14299 9222 16008 9274
rect 1104 9200 16008 9222
rect 4062 9120 4068 9172
rect 4120 9120 4126 9172
rect 4614 9120 4620 9172
rect 4672 9120 4678 9172
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 5537 9163 5595 9169
rect 5537 9160 5549 9163
rect 4856 9132 5549 9160
rect 4856 9120 4862 9132
rect 5537 9129 5549 9132
rect 5583 9129 5595 9163
rect 5537 9123 5595 9129
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8202 9160 8208 9172
rect 8159 9132 8208 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 8202 9120 8208 9132
rect 8260 9160 8266 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 8260 9132 10057 9160
rect 8260 9120 8266 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 11146 9120 11152 9172
rect 11204 9160 11210 9172
rect 14737 9163 14795 9169
rect 11204 9132 12296 9160
rect 11204 9120 11210 9132
rect 2133 9027 2191 9033
rect 2133 8993 2145 9027
rect 2179 9024 2191 9027
rect 4080 9024 4108 9120
rect 12268 9104 12296 9132
rect 12452 9132 13584 9160
rect 12452 9104 12480 9132
rect 5442 9052 5448 9104
rect 5500 9052 5506 9104
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 7248 9064 8524 9092
rect 7248 9052 7254 9064
rect 5460 9024 5488 9052
rect 8202 9024 8208 9036
rect 2179 8996 4108 9024
rect 4356 8996 5488 9024
rect 7116 8996 8208 9024
rect 2179 8993 2191 8996
rect 2133 8987 2191 8993
rect 1854 8916 1860 8968
rect 1912 8916 1918 8968
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 4356 8956 4384 8996
rect 4111 8928 4384 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3252 8820 3280 8916
rect 3108 8792 3280 8820
rect 3605 8823 3663 8829
rect 3108 8780 3114 8792
rect 3605 8789 3617 8823
rect 3651 8820 3663 8823
rect 4080 8820 4108 8919
rect 4522 8916 4528 8968
rect 4580 8956 4586 8968
rect 7116 8965 7144 8996
rect 8202 8984 8208 8996
rect 8260 9024 8266 9036
rect 8260 8996 8432 9024
rect 8260 8984 8266 8996
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4580 8928 4905 8956
rect 4580 8916 4586 8928
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 7248 8928 7297 8956
rect 7248 8916 7254 8928
rect 7285 8925 7297 8928
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 8018 8916 8024 8968
rect 8076 8916 8082 8968
rect 8110 8916 8116 8968
rect 8168 8916 8174 8968
rect 8404 8965 8432 8996
rect 8496 8965 8524 9064
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 8665 9095 8723 9101
rect 8665 9092 8677 9095
rect 8628 9064 8677 9092
rect 8628 9052 8634 9064
rect 8665 9061 8677 9064
rect 8711 9061 8723 9095
rect 8665 9055 8723 9061
rect 11514 9052 11520 9104
rect 11572 9052 11578 9104
rect 11606 9052 11612 9104
rect 11664 9052 11670 9104
rect 12250 9052 12256 9104
rect 12308 9052 12314 9104
rect 12434 9052 12440 9104
rect 12492 9052 12498 9104
rect 13556 9101 13584 9132
rect 14737 9129 14749 9163
rect 14783 9160 14795 9163
rect 15010 9160 15016 9172
rect 14783 9132 15016 9160
rect 14783 9129 14795 9132
rect 14737 9123 14795 9129
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 15378 9120 15384 9172
rect 15436 9160 15442 9172
rect 15473 9163 15531 9169
rect 15473 9160 15485 9163
rect 15436 9132 15485 9160
rect 15436 9120 15442 9132
rect 15473 9129 15485 9132
rect 15519 9129 15531 9163
rect 15473 9123 15531 9129
rect 13449 9095 13507 9101
rect 13449 9092 13461 9095
rect 13096 9064 13461 9092
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 9024 10931 9027
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 10919 8996 10977 9024
rect 10919 8993 10931 8996
rect 10873 8987 10931 8993
rect 10965 8993 10977 8996
rect 11011 8993 11023 9027
rect 10965 8987 11023 8993
rect 11238 8984 11244 9036
rect 11296 8984 11302 9036
rect 11342 9027 11400 9033
rect 11342 8993 11354 9027
rect 11388 9024 11400 9027
rect 11532 9024 11560 9052
rect 11388 8996 11560 9024
rect 11624 9024 11652 9052
rect 13096 9033 13124 9064
rect 13449 9061 13461 9064
rect 13495 9061 13507 9095
rect 13449 9055 13507 9061
rect 13541 9095 13599 9101
rect 13541 9061 13553 9095
rect 13587 9092 13599 9095
rect 13587 9064 15056 9092
rect 13587 9061 13599 9064
rect 13541 9055 13599 9061
rect 13081 9027 13139 9033
rect 13081 9024 13093 9027
rect 11624 8996 13093 9024
rect 11388 8993 11400 8996
rect 11342 8987 11400 8993
rect 13081 8993 13093 8996
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 14458 9024 14464 9036
rect 13311 8996 14464 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 14458 8984 14464 8996
rect 14516 8984 14522 9036
rect 14568 9033 14596 9064
rect 14568 9027 14636 9033
rect 14568 8996 14590 9027
rect 14578 8993 14590 8996
rect 14624 8993 14636 9027
rect 14918 9024 14924 9036
rect 14578 8987 14636 8993
rect 14752 8996 14924 9024
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 8481 8959 8539 8965
rect 8481 8925 8493 8959
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7377 8891 7435 8897
rect 7377 8888 7389 8891
rect 7064 8860 7389 8888
rect 7064 8848 7070 8860
rect 7377 8857 7389 8860
rect 7423 8857 7435 8891
rect 8128 8888 8156 8916
rect 9508 8888 9536 8919
rect 9582 8916 9588 8968
rect 9640 8956 9646 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9640 8928 9873 8956
rect 9640 8916 9646 8928
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8956 10195 8959
rect 10183 8928 10916 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 8128 8860 9536 8888
rect 7377 8851 7435 8857
rect 9766 8848 9772 8900
rect 9824 8888 9830 8900
rect 10152 8888 10180 8919
rect 9824 8860 10180 8888
rect 9824 8848 9830 8860
rect 3651 8792 4108 8820
rect 7285 8823 7343 8829
rect 3651 8789 3663 8792
rect 3605 8783 3663 8789
rect 7285 8789 7297 8823
rect 7331 8820 7343 8823
rect 7926 8820 7932 8832
rect 7331 8792 7932 8820
rect 7331 8789 7343 8792
rect 7285 8783 7343 8789
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 8294 8780 8300 8832
rect 8352 8780 8358 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8812 8792 8953 8820
rect 8812 8780 8818 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 9674 8780 9680 8832
rect 9732 8780 9738 8832
rect 10226 8780 10232 8832
rect 10284 8780 10290 8832
rect 10888 8820 10916 8928
rect 11146 8916 11152 8968
rect 11204 8950 11210 8968
rect 11442 8959 11500 8965
rect 11204 8922 11243 8950
rect 11442 8925 11454 8959
rect 11488 8956 11500 8959
rect 11609 8959 11667 8965
rect 11488 8928 11560 8956
rect 11488 8925 11500 8928
rect 11204 8916 11210 8922
rect 11442 8919 11500 8925
rect 11149 8913 11207 8916
rect 11330 8848 11336 8900
rect 11388 8888 11394 8900
rect 11532 8888 11560 8928
rect 11609 8925 11621 8959
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11388 8860 11560 8888
rect 11388 8848 11394 8860
rect 11624 8820 11652 8919
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 11974 8956 11980 8968
rect 11756 8928 11980 8956
rect 11756 8916 11762 8928
rect 11974 8916 11980 8928
rect 12032 8956 12038 8968
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 12032 8928 12173 8956
rect 12032 8916 12038 8928
rect 12161 8925 12173 8928
rect 12207 8925 12219 8959
rect 12989 8959 13047 8965
rect 12989 8956 13001 8959
rect 12161 8919 12219 8925
rect 12268 8928 13001 8956
rect 11882 8848 11888 8900
rect 11940 8888 11946 8900
rect 12069 8891 12127 8897
rect 12069 8888 12081 8891
rect 11940 8860 12081 8888
rect 11940 8848 11946 8860
rect 12069 8857 12081 8860
rect 12115 8888 12127 8891
rect 12268 8888 12296 8928
rect 12989 8925 13001 8928
rect 13035 8925 13047 8959
rect 12989 8919 13047 8925
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8956 14151 8959
rect 14752 8956 14780 8996
rect 14918 8984 14924 8996
rect 14976 8984 14982 9036
rect 15028 8965 15056 9064
rect 14139 8928 14780 8956
rect 14829 8959 14887 8965
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 14829 8925 14841 8959
rect 14875 8925 14887 8959
rect 14829 8919 14887 8925
rect 15013 8959 15071 8965
rect 15013 8925 15025 8959
rect 15059 8925 15071 8959
rect 15013 8919 15071 8925
rect 12115 8860 12296 8888
rect 12115 8857 12127 8860
rect 12069 8851 12127 8857
rect 12434 8848 12440 8900
rect 12492 8848 12498 8900
rect 12529 8891 12587 8897
rect 12529 8857 12541 8891
rect 12575 8888 12587 8891
rect 13814 8888 13820 8900
rect 12575 8860 13820 8888
rect 12575 8857 12587 8860
rect 12529 8851 12587 8857
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 13909 8891 13967 8897
rect 13909 8857 13921 8891
rect 13955 8888 13967 8891
rect 14461 8891 14519 8897
rect 14461 8888 14473 8891
rect 13955 8860 14473 8888
rect 13955 8857 13967 8860
rect 13909 8851 13967 8857
rect 14292 8832 14320 8860
rect 14461 8857 14473 8860
rect 14507 8857 14519 8891
rect 14844 8888 14872 8919
rect 14461 8851 14519 8857
rect 14752 8860 14872 8888
rect 15565 8891 15623 8897
rect 14752 8832 14780 8860
rect 15565 8857 15577 8891
rect 15611 8888 15623 8891
rect 16022 8888 16028 8900
rect 15611 8860 16028 8888
rect 15611 8857 15623 8860
rect 15565 8851 15623 8857
rect 16022 8848 16028 8860
rect 16080 8848 16086 8900
rect 12158 8820 12164 8832
rect 10888 8792 12164 8820
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12618 8780 12624 8832
rect 12676 8780 12682 8832
rect 14274 8780 14280 8832
rect 14332 8780 14338 8832
rect 14369 8823 14427 8829
rect 14369 8789 14381 8823
rect 14415 8820 14427 8823
rect 14734 8820 14740 8832
rect 14415 8792 14740 8820
rect 14415 8789 14427 8792
rect 14369 8783 14427 8789
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15010 8820 15016 8832
rect 14967 8792 15016 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 1104 8730 16008 8752
rect 1104 8678 3473 8730
rect 3525 8678 3537 8730
rect 3589 8678 3601 8730
rect 3653 8678 3665 8730
rect 3717 8678 3729 8730
rect 3781 8678 7199 8730
rect 7251 8678 7263 8730
rect 7315 8678 7327 8730
rect 7379 8678 7391 8730
rect 7443 8678 7455 8730
rect 7507 8678 10925 8730
rect 10977 8678 10989 8730
rect 11041 8678 11053 8730
rect 11105 8678 11117 8730
rect 11169 8678 11181 8730
rect 11233 8678 14651 8730
rect 14703 8678 14715 8730
rect 14767 8678 14779 8730
rect 14831 8678 14843 8730
rect 14895 8678 14907 8730
rect 14959 8678 16008 8730
rect 1104 8656 16008 8678
rect 4430 8616 4436 8628
rect 2792 8588 4436 8616
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 2792 8489 2820 8588
rect 4430 8576 4436 8588
rect 4488 8576 4494 8628
rect 4522 8576 4528 8628
rect 4580 8576 4586 8628
rect 7282 8616 7288 8628
rect 7024 8588 7288 8616
rect 3050 8508 3056 8560
rect 3108 8548 3114 8560
rect 7024 8548 7052 8588
rect 7282 8576 7288 8588
rect 7340 8616 7346 8628
rect 9401 8619 9459 8625
rect 7340 8588 8340 8616
rect 7340 8576 7346 8588
rect 8312 8557 8340 8588
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 9582 8616 9588 8628
rect 9447 8588 9588 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10226 8616 10232 8628
rect 9876 8588 10232 8616
rect 8297 8551 8355 8557
rect 3108 8520 3542 8548
rect 4724 8520 7130 8548
rect 3108 8508 3114 8520
rect 2777 8483 2835 8489
rect 2777 8480 2789 8483
rect 1912 8452 2789 8480
rect 1912 8440 1918 8452
rect 2777 8449 2789 8452
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8412 3111 8415
rect 4617 8415 4675 8421
rect 4617 8412 4629 8415
rect 3099 8384 4629 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 4617 8381 4629 8384
rect 4663 8381 4675 8415
rect 4617 8375 4675 8381
rect 4724 8344 4752 8520
rect 8297 8517 8309 8551
rect 8343 8517 8355 8551
rect 8297 8511 8355 8517
rect 9125 8551 9183 8557
rect 9125 8517 9137 8551
rect 9171 8548 9183 8551
rect 9214 8548 9220 8560
rect 9171 8520 9220 8548
rect 9171 8517 9183 8520
rect 9125 8511 9183 8517
rect 9214 8508 9220 8520
rect 9272 8508 9278 8560
rect 9766 8548 9772 8560
rect 9508 8520 9772 8548
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 4890 8480 4896 8492
rect 4847 8452 4896 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 4890 8440 4896 8452
rect 4948 8440 4954 8492
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 9508 8489 9536 8520
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 9876 8557 9904 8588
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 12158 8576 12164 8628
rect 12216 8576 12222 8628
rect 12437 8619 12495 8625
rect 12437 8585 12449 8619
rect 12483 8585 12495 8619
rect 12437 8579 12495 8585
rect 9861 8551 9919 8557
rect 9861 8517 9873 8551
rect 9907 8517 9919 8551
rect 12452 8548 12480 8579
rect 14458 8576 14464 8628
rect 14516 8576 14522 8628
rect 12989 8551 13047 8557
rect 12989 8548 13001 8551
rect 12452 8520 13001 8548
rect 9861 8511 9919 8517
rect 12989 8517 13001 8520
rect 13035 8517 13047 8551
rect 12989 8511 13047 8517
rect 13446 8508 13452 8560
rect 13504 8508 13510 8560
rect 15378 8508 15384 8560
rect 15436 8548 15442 8560
rect 15473 8551 15531 8557
rect 15473 8548 15485 8551
rect 15436 8520 15485 8548
rect 15436 8508 15442 8520
rect 15473 8517 15485 8520
rect 15519 8517 15531 8551
rect 15473 8511 15531 8517
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6328 8452 6377 8480
rect 6328 8440 6334 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 6365 8443 6423 8449
rect 8220 8452 9321 8480
rect 5077 8415 5135 8421
rect 5077 8412 5089 8415
rect 4816 8384 5089 8412
rect 4816 8356 4844 8384
rect 5077 8381 5089 8384
rect 5123 8381 5135 8415
rect 5077 8375 5135 8381
rect 6086 8372 6092 8424
rect 6144 8412 6150 8424
rect 6641 8415 6699 8421
rect 6641 8412 6653 8415
rect 6144 8384 6653 8412
rect 6144 8372 6150 8384
rect 6641 8381 6653 8384
rect 6687 8381 6699 8415
rect 6641 8375 6699 8381
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 8220 8412 8248 8452
rect 7156 8384 8248 8412
rect 7156 8372 7162 8384
rect 4080 8316 4752 8344
rect 3234 8236 3240 8288
rect 3292 8276 3298 8288
rect 4080 8276 4108 8316
rect 4798 8304 4804 8356
rect 4856 8304 4862 8356
rect 8864 8344 8892 8452
rect 9309 8449 9321 8452
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 12253 8483 12311 8489
rect 10928 8452 10994 8480
rect 10928 8440 10934 8452
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 12618 8480 12624 8492
rect 12299 8452 12624 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 8938 8372 8944 8424
rect 8996 8412 9002 8424
rect 9585 8415 9643 8421
rect 9585 8412 9597 8415
rect 8996 8384 9597 8412
rect 8996 8372 9002 8384
rect 9585 8381 9597 8384
rect 9631 8381 9643 8415
rect 11054 8412 11060 8424
rect 9585 8375 9643 8381
rect 9692 8384 11060 8412
rect 9692 8344 9720 8384
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 11514 8372 11520 8424
rect 11572 8372 11578 8424
rect 12710 8372 12716 8424
rect 12768 8372 12774 8424
rect 13446 8372 13452 8424
rect 13504 8412 13510 8424
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 13504 8384 14657 8412
rect 13504 8372 13510 8384
rect 14645 8381 14657 8384
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 8864 8316 9720 8344
rect 3292 8248 4108 8276
rect 3292 8236 3298 8248
rect 4982 8236 4988 8288
rect 5040 8236 5046 8288
rect 8110 8236 8116 8288
rect 8168 8236 8174 8288
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 11330 8276 11336 8288
rect 11020 8248 11336 8276
rect 11020 8236 11026 8248
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 1104 8186 16008 8208
rect 1104 8134 2813 8186
rect 2865 8134 2877 8186
rect 2929 8134 2941 8186
rect 2993 8134 3005 8186
rect 3057 8134 3069 8186
rect 3121 8134 6539 8186
rect 6591 8134 6603 8186
rect 6655 8134 6667 8186
rect 6719 8134 6731 8186
rect 6783 8134 6795 8186
rect 6847 8134 10265 8186
rect 10317 8134 10329 8186
rect 10381 8134 10393 8186
rect 10445 8134 10457 8186
rect 10509 8134 10521 8186
rect 10573 8134 13991 8186
rect 14043 8134 14055 8186
rect 14107 8134 14119 8186
rect 14171 8134 14183 8186
rect 14235 8134 14247 8186
rect 14299 8134 16008 8186
rect 1104 8112 16008 8134
rect 3421 8075 3479 8081
rect 3421 8041 3433 8075
rect 3467 8072 3479 8075
rect 3970 8072 3976 8084
rect 3467 8044 3976 8072
rect 3467 8041 3479 8044
rect 3421 8035 3479 8041
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 4709 8075 4767 8081
rect 4709 8072 4721 8075
rect 4488 8044 4721 8072
rect 4488 8032 4494 8044
rect 4709 8041 4721 8044
rect 4755 8041 4767 8075
rect 4709 8035 4767 8041
rect 3605 7939 3663 7945
rect 3605 7905 3617 7939
rect 3651 7936 3663 7939
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 3651 7908 4353 7936
rect 3651 7905 3663 7908
rect 3605 7899 3663 7905
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4724 7936 4752 8035
rect 8018 8032 8024 8084
rect 8076 8072 8082 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 8076 8044 8217 8072
rect 8076 8032 8082 8044
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 8205 8035 8263 8041
rect 8665 8075 8723 8081
rect 8665 8041 8677 8075
rect 8711 8072 8723 8075
rect 8754 8072 8760 8084
rect 8711 8044 8760 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 11514 8072 11520 8084
rect 10735 8044 11520 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 12250 8032 12256 8084
rect 12308 8032 12314 8084
rect 11054 7964 11060 8016
rect 11112 7964 11118 8016
rect 6270 7936 6276 7948
rect 4724 7908 6276 7936
rect 4341 7899 4399 7905
rect 3326 7828 3332 7880
rect 3384 7828 3390 7880
rect 3620 7800 3648 7899
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7936 6607 7939
rect 7006 7936 7012 7948
rect 6595 7908 7012 7936
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 7006 7896 7012 7908
rect 7064 7896 7070 7948
rect 7282 7896 7288 7948
rect 7340 7936 7346 7948
rect 7742 7936 7748 7948
rect 7340 7908 7748 7936
rect 7340 7896 7346 7908
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 7944 7908 8524 7936
rect 7944 7880 7972 7908
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 5442 7868 5448 7880
rect 4203 7840 5448 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 7926 7828 7932 7880
rect 7984 7828 7990 7880
rect 8386 7828 8392 7880
rect 8444 7828 8450 7880
rect 8496 7877 8524 7908
rect 8938 7896 8944 7948
rect 8996 7896 9002 7948
rect 9217 7939 9275 7945
rect 9217 7905 9229 7939
rect 9263 7936 9275 7939
rect 9674 7936 9680 7948
rect 9263 7908 9680 7936
rect 9263 7905 9275 7908
rect 9217 7899 9275 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 12268 7936 12296 8032
rect 13909 8007 13967 8013
rect 13909 7973 13921 8007
rect 13955 8004 13967 8007
rect 14366 8004 14372 8016
rect 13955 7976 14372 8004
rect 13955 7973 13967 7976
rect 13909 7967 13967 7973
rect 14366 7964 14372 7976
rect 14424 8004 14430 8016
rect 14424 7976 15148 8004
rect 14424 7964 14430 7976
rect 15120 7948 15148 7976
rect 11388 7908 12296 7936
rect 12437 7939 12495 7945
rect 11388 7896 11394 7908
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 13814 7936 13820 7948
rect 12483 7908 13820 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 14458 7896 14464 7948
rect 14516 7936 14522 7948
rect 14829 7939 14887 7945
rect 14829 7936 14841 7939
rect 14516 7908 14841 7936
rect 14516 7896 14522 7908
rect 14829 7905 14841 7908
rect 14875 7905 14887 7939
rect 14829 7899 14887 7905
rect 15102 7896 15108 7948
rect 15160 7896 15166 7948
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 10962 7868 10968 7880
rect 10827 7840 10968 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 3344 7772 3648 7800
rect 6181 7803 6239 7809
rect 3344 7744 3372 7772
rect 6181 7769 6193 7803
rect 6227 7769 6239 7803
rect 6181 7763 6239 7769
rect 3326 7692 3332 7744
rect 3384 7692 3390 7744
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 3970 7732 3976 7744
rect 3651 7704 3976 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 4338 7692 4344 7744
rect 4396 7692 4402 7744
rect 6196 7732 6224 7763
rect 6822 7760 6828 7812
rect 6880 7760 6886 7812
rect 7282 7760 7288 7812
rect 7340 7760 7346 7812
rect 8294 7800 8300 7812
rect 8036 7772 8300 7800
rect 6840 7732 6868 7760
rect 6196 7704 6868 7732
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 8036 7741 8064 7772
rect 8294 7760 8300 7772
rect 8352 7800 8358 7812
rect 8772 7800 8800 7831
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7868 11207 7871
rect 11606 7868 11612 7880
rect 11195 7840 11612 7868
rect 11195 7837 11207 7840
rect 11149 7831 11207 7837
rect 11606 7828 11612 7840
rect 11664 7828 11670 7880
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 9214 7800 9220 7812
rect 8352 7772 9220 7800
rect 8352 7760 8358 7772
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 12176 7800 12204 7831
rect 13446 7828 13452 7880
rect 13504 7868 13510 7880
rect 14737 7871 14795 7877
rect 13504 7840 13570 7868
rect 13504 7828 13510 7840
rect 14737 7837 14749 7871
rect 14783 7868 14795 7871
rect 15194 7868 15200 7880
rect 14783 7840 15200 7868
rect 14783 7837 14795 7840
rect 14737 7831 14795 7837
rect 15194 7828 15200 7840
rect 15252 7828 15258 7880
rect 12710 7800 12716 7812
rect 10442 7772 10824 7800
rect 12176 7772 12716 7800
rect 10796 7744 10824 7772
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 6972 7704 8033 7732
rect 6972 7692 6978 7704
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 10778 7692 10784 7744
rect 10836 7692 10842 7744
rect 14093 7735 14151 7741
rect 14093 7701 14105 7735
rect 14139 7732 14151 7735
rect 14366 7732 14372 7744
rect 14139 7704 14372 7732
rect 14139 7701 14151 7704
rect 14093 7695 14151 7701
rect 14366 7692 14372 7704
rect 14424 7692 14430 7744
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 15344 7704 15485 7732
rect 15344 7692 15350 7704
rect 15473 7701 15485 7704
rect 15519 7701 15531 7735
rect 15473 7695 15531 7701
rect 1104 7642 16008 7664
rect 1104 7590 3473 7642
rect 3525 7590 3537 7642
rect 3589 7590 3601 7642
rect 3653 7590 3665 7642
rect 3717 7590 3729 7642
rect 3781 7590 7199 7642
rect 7251 7590 7263 7642
rect 7315 7590 7327 7642
rect 7379 7590 7391 7642
rect 7443 7590 7455 7642
rect 7507 7590 10925 7642
rect 10977 7590 10989 7642
rect 11041 7590 11053 7642
rect 11105 7590 11117 7642
rect 11169 7590 11181 7642
rect 11233 7590 14651 7642
rect 14703 7590 14715 7642
rect 14767 7590 14779 7642
rect 14831 7590 14843 7642
rect 14895 7590 14907 7642
rect 14959 7590 16008 7642
rect 1104 7568 16008 7590
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 3292 7500 3556 7528
rect 3292 7488 3298 7500
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 1912 7364 2145 7392
rect 1912 7352 1918 7364
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 3528 7378 3556 7500
rect 4246 7488 4252 7540
rect 4304 7488 4310 7540
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 4396 7500 4445 7528
rect 4396 7488 4402 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 4433 7491 4491 7497
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 5500 7500 5733 7528
rect 5500 7488 5506 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 5721 7491 5779 7497
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6052 7500 8156 7528
rect 6052 7488 6058 7500
rect 4264 7460 4292 7488
rect 5261 7463 5319 7469
rect 4264 7432 4568 7460
rect 2133 7355 2191 7361
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 3936 7364 4077 7392
rect 3936 7352 3942 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4338 7352 4344 7404
rect 4396 7352 4402 7404
rect 4540 7401 4568 7432
rect 5261 7429 5273 7463
rect 5307 7460 5319 7463
rect 7006 7460 7012 7472
rect 5307 7432 7012 7460
rect 5307 7429 5319 7432
rect 5261 7423 5319 7429
rect 7006 7420 7012 7432
rect 7064 7420 7070 7472
rect 7742 7420 7748 7472
rect 7800 7420 7806 7472
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 5074 7352 5080 7404
rect 5132 7352 5138 7404
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 5276 7364 5365 7392
rect 5276 7336 5304 7364
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5353 7355 5411 7361
rect 5460 7364 5825 7392
rect 2409 7327 2467 7333
rect 2409 7293 2421 7327
rect 2455 7324 2467 7327
rect 2455 7296 4016 7324
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 3988 7256 4016 7296
rect 4154 7284 4160 7336
rect 4212 7284 4218 7336
rect 4982 7284 4988 7336
rect 5040 7284 5046 7336
rect 5258 7284 5264 7336
rect 5316 7284 5322 7336
rect 4890 7256 4896 7268
rect 3988 7228 4896 7256
rect 4890 7216 4896 7228
rect 4948 7216 4954 7268
rect 5000 7256 5028 7284
rect 5077 7259 5135 7265
rect 5077 7256 5089 7259
rect 5000 7228 5089 7256
rect 5077 7225 5089 7228
rect 5123 7256 5135 7259
rect 5460 7256 5488 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6457 7395 6515 7401
rect 6457 7392 6469 7395
rect 6328 7364 6469 7392
rect 6328 7352 6334 7364
rect 6457 7361 6469 7364
rect 6503 7361 6515 7395
rect 6457 7355 6515 7361
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7324 6791 7327
rect 7190 7324 7196 7336
rect 6779 7296 7196 7324
rect 6779 7293 6791 7296
rect 6733 7287 6791 7293
rect 5123 7228 5488 7256
rect 5644 7256 5672 7287
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 8128 7256 8156 7500
rect 8202 7488 8208 7540
rect 8260 7488 8266 7540
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 9677 7531 9735 7537
rect 9677 7528 9689 7531
rect 8444 7500 9689 7528
rect 8444 7488 8450 7500
rect 9677 7497 9689 7500
rect 9723 7497 9735 7531
rect 9677 7491 9735 7497
rect 11330 7488 11336 7540
rect 11388 7528 11394 7540
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 11388 7500 11621 7528
rect 11388 7488 11394 7500
rect 11609 7497 11621 7500
rect 11655 7497 11667 7531
rect 11609 7491 11667 7497
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 12768 7500 14780 7528
rect 12768 7488 12774 7500
rect 8220 7392 8248 7488
rect 8570 7420 8576 7472
rect 8628 7460 8634 7472
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 8628 7432 9505 7460
rect 8628 7420 8634 7432
rect 9493 7429 9505 7432
rect 9539 7460 9551 7463
rect 9539 7432 9720 7460
rect 9539 7429 9551 7432
rect 9493 7423 9551 7429
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 8220 7364 8953 7392
rect 8941 7361 8953 7364
rect 8987 7392 8999 7395
rect 9125 7395 9183 7401
rect 9125 7392 9137 7395
rect 8987 7364 9137 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9125 7361 9137 7364
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9692 7401 9720 7432
rect 13446 7420 13452 7472
rect 13504 7420 13510 7472
rect 14366 7420 14372 7472
rect 14424 7460 14430 7472
rect 14461 7463 14519 7469
rect 14461 7460 14473 7463
rect 14424 7432 14473 7460
rect 14424 7420 14430 7432
rect 14461 7429 14473 7432
rect 14507 7429 14519 7463
rect 14461 7423 14519 7429
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9272 7364 9597 7392
rect 9272 7352 9278 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9600 7324 9628 7355
rect 9876 7324 9904 7355
rect 11698 7352 11704 7404
rect 11756 7352 11762 7404
rect 14752 7401 14780 7500
rect 15102 7488 15108 7540
rect 15160 7528 15166 7540
rect 15160 7500 15516 7528
rect 15160 7488 15166 7500
rect 14829 7463 14887 7469
rect 14829 7429 14841 7463
rect 14875 7460 14887 7463
rect 15194 7460 15200 7472
rect 14875 7432 15200 7460
rect 14875 7429 14887 7432
rect 14829 7423 14887 7429
rect 15194 7420 15200 7432
rect 15252 7420 15258 7472
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 15010 7352 15016 7404
rect 15068 7352 15074 7404
rect 15102 7352 15108 7404
rect 15160 7352 15166 7404
rect 15488 7401 15516 7500
rect 15381 7395 15439 7401
rect 15381 7392 15393 7395
rect 15212 7364 15393 7392
rect 9600 7296 9904 7324
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 12989 7327 13047 7333
rect 12989 7324 13001 7327
rect 12492 7296 13001 7324
rect 12492 7284 12498 7296
rect 12989 7293 13001 7296
rect 13035 7324 13047 7327
rect 14918 7324 14924 7336
rect 13035 7296 14924 7324
rect 13035 7293 13047 7296
rect 12989 7287 13047 7293
rect 14918 7284 14924 7296
rect 14976 7324 14982 7336
rect 15212 7324 15240 7364
rect 15381 7361 15393 7364
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 14976 7296 15240 7324
rect 14976 7284 14982 7296
rect 15286 7284 15292 7336
rect 15344 7284 15350 7336
rect 9674 7256 9680 7268
rect 5644 7228 6592 7256
rect 8128 7228 9680 7256
rect 5123 7225 5135 7228
rect 5077 7219 5135 7225
rect 3418 7148 3424 7200
rect 3476 7188 3482 7200
rect 3881 7191 3939 7197
rect 3881 7188 3893 7191
rect 3476 7160 3893 7188
rect 3476 7148 3482 7160
rect 3881 7157 3893 7160
rect 3927 7188 3939 7191
rect 4246 7188 4252 7200
rect 3927 7160 4252 7188
rect 3927 7157 3939 7160
rect 3881 7151 3939 7157
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 4801 7191 4859 7197
rect 4801 7157 4813 7191
rect 4847 7188 4859 7191
rect 5994 7188 6000 7200
rect 4847 7160 6000 7188
rect 4847 7157 4859 7160
rect 4801 7151 4859 7157
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6178 7148 6184 7200
rect 6236 7148 6242 7200
rect 6564 7188 6592 7228
rect 9674 7216 9680 7228
rect 9732 7216 9738 7268
rect 15102 7216 15108 7268
rect 15160 7256 15166 7268
rect 15565 7259 15623 7265
rect 15565 7256 15577 7259
rect 15160 7228 15577 7256
rect 15160 7216 15166 7228
rect 15565 7225 15577 7228
rect 15611 7225 15623 7259
rect 15565 7219 15623 7225
rect 8110 7188 8116 7200
rect 6564 7160 8116 7188
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8386 7148 8392 7200
rect 8444 7148 8450 7200
rect 9306 7148 9312 7200
rect 9364 7148 9370 7200
rect 1104 7098 16008 7120
rect 1104 7046 2813 7098
rect 2865 7046 2877 7098
rect 2929 7046 2941 7098
rect 2993 7046 3005 7098
rect 3057 7046 3069 7098
rect 3121 7046 6539 7098
rect 6591 7046 6603 7098
rect 6655 7046 6667 7098
rect 6719 7046 6731 7098
rect 6783 7046 6795 7098
rect 6847 7046 10265 7098
rect 10317 7046 10329 7098
rect 10381 7046 10393 7098
rect 10445 7046 10457 7098
rect 10509 7046 10521 7098
rect 10573 7046 13991 7098
rect 14043 7046 14055 7098
rect 14107 7046 14119 7098
rect 14171 7046 14183 7098
rect 14235 7046 14247 7098
rect 14299 7046 16008 7098
rect 1104 7024 16008 7046
rect 2120 6987 2178 6993
rect 2120 6953 2132 6987
rect 2166 6984 2178 6987
rect 4154 6984 4160 6996
rect 2166 6956 4160 6984
rect 2166 6953 2178 6956
rect 2120 6947 2178 6953
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 4890 6944 4896 6996
rect 4948 6944 4954 6996
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5629 6987 5687 6993
rect 5629 6984 5641 6987
rect 5132 6956 5641 6984
rect 5132 6944 5138 6956
rect 5629 6953 5641 6956
rect 5675 6953 5687 6987
rect 5629 6947 5687 6953
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 7248 6956 7573 6984
rect 7248 6944 7254 6956
rect 7561 6953 7573 6956
rect 7607 6953 7619 6987
rect 7561 6947 7619 6953
rect 8202 6944 8208 6996
rect 8260 6944 8266 6996
rect 10492 6987 10550 6993
rect 10492 6953 10504 6987
rect 10538 6984 10550 6987
rect 11514 6984 11520 6996
rect 10538 6956 11520 6984
rect 10538 6953 10550 6956
rect 10492 6947 10550 6953
rect 11514 6944 11520 6956
rect 11572 6944 11578 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 11977 6987 12035 6993
rect 11977 6984 11989 6987
rect 11756 6956 11989 6984
rect 11756 6944 11762 6956
rect 11977 6953 11989 6956
rect 12023 6953 12035 6987
rect 11977 6947 12035 6953
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13872 6956 14105 6984
rect 13872 6944 13878 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 3973 6919 4031 6925
rect 3973 6885 3985 6919
rect 4019 6916 4031 6919
rect 4062 6916 4068 6928
rect 4019 6888 4068 6916
rect 4019 6885 4031 6888
rect 3973 6879 4031 6885
rect 4062 6876 4068 6888
rect 4120 6876 4126 6928
rect 5258 6876 5264 6928
rect 5316 6916 5322 6928
rect 6730 6916 6736 6928
rect 5316 6888 6736 6916
rect 5316 6876 5322 6888
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 8220 6916 8248 6944
rect 12710 6916 12716 6928
rect 7392 6888 8248 6916
rect 12406 6888 12716 6916
rect 1854 6808 1860 6860
rect 1912 6808 1918 6860
rect 4080 6848 4108 6876
rect 4801 6851 4859 6857
rect 4080 6820 4384 6848
rect 3234 6740 3240 6792
rect 3292 6740 3298 6792
rect 4065 6783 4123 6789
rect 4065 6780 4077 6783
rect 3988 6752 4077 6780
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3252 6644 3280 6740
rect 3988 6656 4016 6752
rect 4065 6749 4077 6752
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4246 6780 4252 6792
rect 4203 6752 4252 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 3108 6616 3280 6644
rect 3605 6647 3663 6653
rect 3108 6604 3114 6616
rect 3605 6613 3617 6647
rect 3651 6644 3663 6647
rect 3970 6644 3976 6656
rect 3651 6616 3976 6644
rect 3651 6613 3663 6616
rect 3605 6607 3663 6613
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4172 6644 4200 6743
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4356 6780 4384 6820
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 4847 6820 5365 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 7009 6851 7067 6857
rect 7009 6848 7021 6851
rect 5500 6820 7021 6848
rect 5500 6808 5506 6820
rect 7009 6817 7021 6820
rect 7055 6817 7067 6851
rect 7009 6811 7067 6817
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 7392 6857 7420 6888
rect 7377 6851 7435 6857
rect 7377 6848 7389 6851
rect 7156 6820 7389 6848
rect 7156 6808 7162 6820
rect 7377 6817 7389 6820
rect 7423 6817 7435 6851
rect 7926 6848 7932 6860
rect 7377 6811 7435 6817
rect 7668 6820 7932 6848
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4356 6752 5089 6780
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5166 6740 5172 6792
rect 5224 6740 5230 6792
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 5460 6780 5488 6808
rect 5307 6752 5488 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 5626 6740 5632 6792
rect 5684 6740 5690 6792
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 6178 6780 6184 6792
rect 6043 6752 6184 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6730 6740 6736 6792
rect 6788 6740 6794 6792
rect 7282 6740 7288 6792
rect 7340 6740 7346 6792
rect 7668 6780 7696 6820
rect 7852 6789 7880 6820
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8570 6848 8576 6860
rect 8067 6820 8576 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 10229 6851 10287 6857
rect 10229 6817 10241 6851
rect 10275 6848 10287 6851
rect 12406 6848 12434 6888
rect 12710 6876 12716 6888
rect 12768 6876 12774 6928
rect 14737 6919 14795 6925
rect 14737 6885 14749 6919
rect 14783 6885 14795 6919
rect 14737 6879 14795 6885
rect 14366 6848 14372 6860
rect 10275 6820 12434 6848
rect 14292 6820 14372 6848
rect 10275 6817 10287 6820
rect 10229 6811 10287 6817
rect 7392 6752 7696 6780
rect 7745 6783 7803 6789
rect 4430 6672 4436 6724
rect 4488 6712 4494 6724
rect 5721 6715 5779 6721
rect 5721 6712 5733 6715
rect 4488 6684 5733 6712
rect 4488 6672 4494 6684
rect 5721 6681 5733 6684
rect 5767 6681 5779 6715
rect 5721 6675 5779 6681
rect 5905 6715 5963 6721
rect 5905 6681 5917 6715
rect 5951 6681 5963 6715
rect 5905 6675 5963 6681
rect 5920 6644 5948 6675
rect 6086 6672 6092 6724
rect 6144 6672 6150 6724
rect 7006 6672 7012 6724
rect 7064 6712 7070 6724
rect 7392 6712 7420 6752
rect 7745 6749 7757 6783
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8386 6780 8392 6792
rect 8159 6752 8392 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 7064 6684 7420 6712
rect 7760 6712 7788 6743
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 12066 6740 12072 6792
rect 12124 6780 12130 6792
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12124 6752 12725 6780
rect 12124 6740 12130 6752
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 13906 6740 13912 6792
rect 13964 6740 13970 6792
rect 14292 6789 14320 6820
rect 14366 6808 14372 6820
rect 14424 6848 14430 6860
rect 14752 6848 14780 6879
rect 14424 6820 14780 6848
rect 14424 6808 14430 6820
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14458 6740 14464 6792
rect 14516 6780 14522 6792
rect 14553 6783 14611 6789
rect 14553 6780 14565 6783
rect 14516 6752 14565 6780
rect 14516 6740 14522 6752
rect 14553 6749 14565 6752
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 14918 6740 14924 6792
rect 14976 6780 14982 6792
rect 15013 6783 15071 6789
rect 15013 6780 15025 6783
rect 14976 6752 15025 6780
rect 14976 6740 14982 6752
rect 15013 6749 15025 6752
rect 15059 6749 15071 6783
rect 15013 6743 15071 6749
rect 8294 6712 8300 6724
rect 7760 6684 8300 6712
rect 7064 6672 7070 6684
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 10778 6672 10784 6724
rect 10836 6712 10842 6724
rect 13446 6712 13452 6724
rect 10836 6684 10994 6712
rect 11808 6684 13452 6712
rect 10836 6672 10842 6684
rect 4172 6616 5948 6644
rect 6104 6644 6132 6672
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 6104 6616 6193 6644
rect 6181 6613 6193 6616
rect 6227 6613 6239 6647
rect 10888 6644 10916 6684
rect 11808 6644 11836 6684
rect 13446 6672 13452 6684
rect 13504 6672 13510 6724
rect 10888 6616 11836 6644
rect 6181 6607 6239 6613
rect 12158 6604 12164 6656
rect 12216 6604 12222 6656
rect 13924 6644 13952 6740
rect 14737 6715 14795 6721
rect 14737 6712 14749 6715
rect 14476 6684 14749 6712
rect 14476 6653 14504 6684
rect 14737 6681 14749 6684
rect 14783 6712 14795 6715
rect 15102 6712 15108 6724
rect 14783 6684 15108 6712
rect 14783 6681 14795 6684
rect 14737 6675 14795 6681
rect 15102 6672 15108 6684
rect 15160 6672 15166 6724
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 13924 6616 14473 6644
rect 14461 6613 14473 6616
rect 14507 6613 14519 6647
rect 14461 6607 14519 6613
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 14608 6616 14933 6644
rect 14608 6604 14614 6616
rect 14921 6613 14933 6616
rect 14967 6613 14979 6647
rect 14921 6607 14979 6613
rect 1104 6554 16008 6576
rect 1104 6502 3473 6554
rect 3525 6502 3537 6554
rect 3589 6502 3601 6554
rect 3653 6502 3665 6554
rect 3717 6502 3729 6554
rect 3781 6502 7199 6554
rect 7251 6502 7263 6554
rect 7315 6502 7327 6554
rect 7379 6502 7391 6554
rect 7443 6502 7455 6554
rect 7507 6502 10925 6554
rect 10977 6502 10989 6554
rect 11041 6502 11053 6554
rect 11105 6502 11117 6554
rect 11169 6502 11181 6554
rect 11233 6502 14651 6554
rect 14703 6502 14715 6554
rect 14767 6502 14779 6554
rect 14831 6502 14843 6554
rect 14895 6502 14907 6554
rect 14959 6502 16008 6554
rect 1104 6480 16008 6502
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 3252 6412 3433 6440
rect 3252 6384 3280 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 3421 6403 3479 6409
rect 3878 6400 3884 6452
rect 3936 6400 3942 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 5169 6443 5227 6449
rect 5169 6440 5181 6443
rect 4212 6412 5181 6440
rect 4212 6400 4218 6412
rect 5169 6409 5181 6412
rect 5215 6409 5227 6443
rect 5169 6403 5227 6409
rect 7098 6400 7104 6452
rect 7156 6400 7162 6452
rect 8294 6400 8300 6452
rect 8352 6400 8358 6452
rect 11514 6400 11520 6452
rect 11572 6400 11578 6452
rect 12158 6400 12164 6452
rect 12216 6400 12222 6452
rect 3234 6332 3240 6384
rect 3292 6332 3298 6384
rect 3896 6372 3924 6400
rect 3896 6344 5212 6372
rect 5184 6316 5212 6344
rect 3142 6264 3148 6316
rect 3200 6264 3206 6316
rect 3326 6264 3332 6316
rect 3384 6264 3390 6316
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6304 3847 6307
rect 4062 6304 4068 6316
rect 3835 6276 4068 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 3160 6168 3188 6264
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6236 3295 6239
rect 3344 6236 3372 6264
rect 3283 6208 3372 6236
rect 3283 6205 3295 6208
rect 3237 6199 3295 6205
rect 3436 6168 3464 6267
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4430 6264 4436 6316
rect 4488 6264 4494 6316
rect 4614 6264 4620 6316
rect 4672 6264 4678 6316
rect 4893 6307 4951 6313
rect 4893 6273 4905 6307
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5074 6304 5080 6316
rect 5031 6276 5080 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 4448 6236 4476 6264
rect 4028 6208 4476 6236
rect 4908 6236 4936 6267
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5166 6264 5172 6316
rect 5224 6264 5230 6316
rect 5442 6264 5448 6316
rect 5500 6264 5506 6316
rect 7116 6304 7144 6400
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 7116 6276 7205 6304
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 7193 6267 7251 6273
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6304 7435 6307
rect 8312 6304 8340 6400
rect 12176 6372 12204 6400
rect 11992 6344 12204 6372
rect 7423 6276 8340 6304
rect 7423 6273 7435 6276
rect 7377 6267 7435 6273
rect 8938 6264 8944 6316
rect 8996 6304 9002 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 8996 6276 9597 6304
rect 8996 6264 9002 6276
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 10870 6264 10876 6316
rect 10928 6304 10934 6316
rect 11701 6307 11759 6313
rect 10928 6276 10994 6304
rect 10928 6264 10934 6276
rect 11701 6273 11713 6307
rect 11747 6304 11759 6307
rect 11882 6304 11888 6316
rect 11747 6276 11888 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 11992 6313 12020 6344
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 12066 6264 12072 6316
rect 12124 6264 12130 6316
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 5460 6236 5488 6264
rect 4908 6208 5488 6236
rect 4028 6196 4034 6208
rect 9858 6196 9864 6248
rect 9916 6196 9922 6248
rect 11333 6239 11391 6245
rect 11333 6205 11345 6239
rect 11379 6236 11391 6239
rect 12084 6236 12112 6264
rect 11379 6208 12112 6236
rect 11379 6205 11391 6208
rect 11333 6199 11391 6205
rect 5626 6168 5632 6180
rect 3160 6140 5632 6168
rect 5626 6128 5632 6140
rect 5684 6128 5690 6180
rect 11698 6128 11704 6180
rect 11756 6168 11762 6180
rect 12176 6168 12204 6267
rect 12342 6168 12348 6180
rect 11756 6140 12348 6168
rect 11756 6128 11762 6140
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 4709 6103 4767 6109
rect 4709 6100 4721 6103
rect 4571 6072 4721 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 4709 6069 4721 6072
rect 4755 6069 4767 6103
rect 4709 6063 4767 6069
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 7285 6103 7343 6109
rect 7285 6100 7297 6103
rect 7156 6072 7297 6100
rect 7156 6060 7162 6072
rect 7285 6069 7297 6072
rect 7331 6069 7343 6103
rect 7285 6063 7343 6069
rect 1104 6010 16008 6032
rect 1104 5958 2813 6010
rect 2865 5958 2877 6010
rect 2929 5958 2941 6010
rect 2993 5958 3005 6010
rect 3057 5958 3069 6010
rect 3121 5958 6539 6010
rect 6591 5958 6603 6010
rect 6655 5958 6667 6010
rect 6719 5958 6731 6010
rect 6783 5958 6795 6010
rect 6847 5958 10265 6010
rect 10317 5958 10329 6010
rect 10381 5958 10393 6010
rect 10445 5958 10457 6010
rect 10509 5958 10521 6010
rect 10573 5958 13991 6010
rect 14043 5958 14055 6010
rect 14107 5958 14119 6010
rect 14171 5958 14183 6010
rect 14235 5958 14247 6010
rect 14299 5958 16008 6010
rect 1104 5936 16008 5958
rect 4430 5896 4436 5908
rect 3160 5868 4436 5896
rect 3160 5837 3188 5868
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 9858 5856 9864 5908
rect 9916 5896 9922 5908
rect 10137 5899 10195 5905
rect 10137 5896 10149 5899
rect 9916 5868 10149 5896
rect 9916 5856 9922 5868
rect 10137 5865 10149 5868
rect 10183 5865 10195 5899
rect 10137 5859 10195 5865
rect 3145 5831 3203 5837
rect 3145 5797 3157 5831
rect 3191 5797 3203 5831
rect 3145 5791 3203 5797
rect 4065 5831 4123 5837
rect 4065 5797 4077 5831
rect 4111 5828 4123 5831
rect 4706 5828 4712 5840
rect 4111 5800 4712 5828
rect 4111 5797 4123 5800
rect 4065 5791 4123 5797
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 12529 5831 12587 5837
rect 12529 5797 12541 5831
rect 12575 5828 12587 5831
rect 12618 5828 12624 5840
rect 12575 5800 12624 5828
rect 12575 5797 12587 5800
rect 12529 5791 12587 5797
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 14366 5788 14372 5840
rect 14424 5828 14430 5840
rect 14424 5800 14688 5828
rect 14424 5788 14430 5800
rect 5534 5760 5540 5772
rect 2700 5732 5540 5760
rect 2700 5704 2728 5732
rect 2682 5652 2688 5704
rect 2740 5652 2746 5704
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 3068 5624 3096 5655
rect 3234 5652 3240 5704
rect 3292 5652 3298 5704
rect 3326 5652 3332 5704
rect 3384 5652 3390 5704
rect 3528 5701 3556 5732
rect 5534 5720 5540 5732
rect 5592 5720 5598 5772
rect 6917 5763 6975 5769
rect 6917 5729 6929 5763
rect 6963 5729 6975 5763
rect 12894 5760 12900 5772
rect 6917 5723 6975 5729
rect 12268 5732 12900 5760
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5661 3571 5695
rect 3513 5655 3571 5661
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 3970 5692 3976 5704
rect 3835 5664 3976 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 6454 5692 6460 5704
rect 6196 5664 6460 5692
rect 2832 5596 3280 5624
rect 2832 5584 2838 5596
rect 2869 5559 2927 5565
rect 2869 5525 2881 5559
rect 2915 5556 2927 5559
rect 3142 5556 3148 5568
rect 2915 5528 3148 5556
rect 2915 5525 2927 5528
rect 2869 5519 2927 5525
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 3252 5556 3280 5596
rect 3878 5584 3884 5636
rect 3936 5584 3942 5636
rect 4062 5584 4068 5636
rect 4120 5584 4126 5636
rect 4080 5556 4108 5584
rect 6196 5568 6224 5664
rect 6454 5652 6460 5664
rect 6512 5692 6518 5704
rect 6733 5695 6791 5701
rect 6733 5692 6745 5695
rect 6512 5664 6745 5692
rect 6512 5652 6518 5664
rect 6733 5661 6745 5664
rect 6779 5661 6791 5695
rect 6932 5692 6960 5723
rect 7006 5692 7012 5704
rect 6932 5664 7012 5692
rect 6733 5655 6791 5661
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 10321 5695 10379 5701
rect 7147 5664 8616 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 8588 5568 8616 5664
rect 10321 5661 10333 5695
rect 10367 5661 10379 5695
rect 10321 5655 10379 5661
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10594 5692 10600 5704
rect 10459 5664 10600 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 10336 5624 10364 5655
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12268 5701 12296 5732
rect 12894 5720 12900 5732
rect 12952 5720 12958 5772
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5760 14151 5763
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14139 5732 14565 5760
rect 14139 5729 14151 5732
rect 14093 5723 14151 5729
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 12253 5695 12311 5701
rect 12253 5692 12265 5695
rect 12032 5664 12265 5692
rect 12032 5652 12038 5664
rect 12253 5661 12265 5664
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 12342 5652 12348 5704
rect 12400 5652 12406 5704
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13964 5664 14289 5692
rect 13964 5652 13970 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 14458 5692 14464 5704
rect 14415 5664 14464 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 14660 5701 14688 5800
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 15378 5652 15384 5704
rect 15436 5652 15442 5704
rect 11514 5624 11520 5636
rect 10336 5596 11520 5624
rect 11514 5584 11520 5596
rect 11572 5584 11578 5636
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 12529 5627 12587 5633
rect 12529 5624 12541 5627
rect 12492 5596 12541 5624
rect 12492 5584 12498 5596
rect 12529 5593 12541 5596
rect 12575 5593 12587 5627
rect 14476 5624 14504 5652
rect 14829 5627 14887 5633
rect 14829 5624 14841 5627
rect 14476 5596 14841 5624
rect 12529 5587 12587 5593
rect 14829 5593 14841 5596
rect 14875 5593 14887 5627
rect 14829 5587 14887 5593
rect 3252 5528 4108 5556
rect 6178 5516 6184 5568
rect 6236 5516 6242 5568
rect 6822 5516 6828 5568
rect 6880 5516 6886 5568
rect 7009 5559 7067 5565
rect 7009 5525 7021 5559
rect 7055 5556 7067 5559
rect 8294 5556 8300 5568
rect 7055 5528 8300 5556
rect 7055 5525 7067 5528
rect 7009 5519 7067 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8570 5516 8576 5568
rect 8628 5516 8634 5568
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 11701 5559 11759 5565
rect 11701 5556 11713 5559
rect 8996 5528 11713 5556
rect 8996 5516 9002 5528
rect 11701 5525 11713 5528
rect 11747 5556 11759 5559
rect 12710 5556 12716 5568
rect 11747 5528 12716 5556
rect 11747 5525 11759 5528
rect 11701 5519 11759 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 14090 5516 14096 5568
rect 14148 5516 14154 5568
rect 1104 5466 16008 5488
rect 1104 5414 3473 5466
rect 3525 5414 3537 5466
rect 3589 5414 3601 5466
rect 3653 5414 3665 5466
rect 3717 5414 3729 5466
rect 3781 5414 7199 5466
rect 7251 5414 7263 5466
rect 7315 5414 7327 5466
rect 7379 5414 7391 5466
rect 7443 5414 7455 5466
rect 7507 5414 10925 5466
rect 10977 5414 10989 5466
rect 11041 5414 11053 5466
rect 11105 5414 11117 5466
rect 11169 5414 11181 5466
rect 11233 5414 14651 5466
rect 14703 5414 14715 5466
rect 14767 5414 14779 5466
rect 14831 5414 14843 5466
rect 14895 5414 14907 5466
rect 14959 5414 16008 5466
rect 1104 5392 16008 5414
rect 3053 5355 3111 5361
rect 3053 5321 3065 5355
rect 3099 5352 3111 5355
rect 3326 5352 3332 5364
rect 3099 5324 3332 5352
rect 3099 5321 3111 5324
rect 3053 5315 3111 5321
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 4614 5352 4620 5364
rect 4479 5324 4620 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 3970 5284 3976 5296
rect 2976 5256 3976 5284
rect 2976 5225 3004 5256
rect 3970 5244 3976 5256
rect 4028 5284 4034 5296
rect 4448 5284 4476 5315
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 7616 5324 9674 5352
rect 7616 5312 7622 5324
rect 4028 5256 4476 5284
rect 4028 5244 4034 5256
rect 6086 5244 6092 5296
rect 6144 5284 6150 5296
rect 6144 5256 7696 5284
rect 6144 5244 6150 5256
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3418 5216 3424 5228
rect 3108 5188 3424 5216
rect 3108 5176 3114 5188
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5216 3755 5219
rect 3878 5216 3884 5228
rect 3743 5188 3884 5216
rect 3743 5185 3755 5188
rect 3697 5179 3755 5185
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5216 4767 5219
rect 4982 5216 4988 5228
rect 4755 5188 4988 5216
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 6178 5176 6184 5228
rect 6236 5176 6242 5228
rect 6380 5225 6408 5256
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5216 6975 5219
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 6963 5188 7389 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5148 2743 5151
rect 3326 5148 3332 5160
rect 2731 5120 3332 5148
rect 2731 5117 2743 5120
rect 2685 5111 2743 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3786 5108 3792 5160
rect 3844 5108 3850 5160
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4890 5148 4896 5160
rect 4120 5120 4896 5148
rect 4120 5108 4126 5120
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 6748 5148 6776 5179
rect 7392 5148 7420 5179
rect 7558 5176 7564 5228
rect 7616 5176 7622 5228
rect 7668 5225 7696 5256
rect 7760 5256 9352 5284
rect 7760 5225 7788 5256
rect 9324 5228 9352 5256
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 7929 5181 7987 5187
rect 7929 5178 7941 5181
rect 7852 5150 7941 5178
rect 7852 5148 7880 5150
rect 6748 5120 7328 5148
rect 7392 5120 7880 5148
rect 7929 5147 7941 5150
rect 7975 5147 7987 5181
rect 9306 5176 9312 5228
rect 9364 5176 9370 5228
rect 7929 5141 7987 5147
rect 2869 5083 2927 5089
rect 2869 5049 2881 5083
rect 2915 5080 2927 5083
rect 5166 5080 5172 5092
rect 2915 5052 5172 5080
rect 2915 5049 2927 5052
rect 2869 5043 2927 5049
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 5442 5040 5448 5092
rect 5500 5080 5506 5092
rect 6457 5083 6515 5089
rect 6457 5080 6469 5083
rect 5500 5052 6469 5080
rect 5500 5040 5506 5052
rect 6457 5049 6469 5052
rect 6503 5049 6515 5083
rect 6457 5043 6515 5049
rect 2498 4972 2504 5024
rect 2556 5012 2562 5024
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 2556 4984 2789 5012
rect 2556 4972 2562 4984
rect 2777 4981 2789 4984
rect 2823 4981 2835 5015
rect 2777 4975 2835 4981
rect 3234 4972 3240 5024
rect 3292 5012 3298 5024
rect 4062 5012 4068 5024
rect 3292 4984 4068 5012
rect 3292 4972 3298 4984
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4614 4972 4620 5024
rect 4672 4972 4678 5024
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 6822 5012 6828 5024
rect 6052 4984 6828 5012
rect 6052 4972 6058 4984
rect 6822 4972 6828 4984
rect 6880 5012 6886 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6880 4984 7205 5012
rect 6880 4972 6886 4984
rect 7193 4981 7205 4984
rect 7239 4981 7251 5015
rect 7300 5012 7328 5120
rect 7668 5092 7696 5120
rect 7650 5040 7656 5092
rect 7708 5040 7714 5092
rect 7558 5012 7564 5024
rect 7300 4984 7564 5012
rect 7193 4975 7251 4981
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 7837 5015 7895 5021
rect 7837 4981 7849 5015
rect 7883 5012 7895 5015
rect 9122 5012 9128 5024
rect 7883 4984 9128 5012
rect 7883 4981 7895 4984
rect 7837 4975 7895 4981
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9214 4972 9220 5024
rect 9272 4972 9278 5024
rect 9646 5012 9674 5324
rect 11514 5312 11520 5364
rect 11572 5312 11578 5364
rect 11885 5355 11943 5361
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 11931 5324 12664 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 12342 5244 12348 5296
rect 12400 5284 12406 5296
rect 12400 5256 12572 5284
rect 12400 5244 12406 5256
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10594 5216 10600 5228
rect 10091 5188 10600 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 10594 5176 10600 5188
rect 10652 5216 10658 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10652 5188 10977 5216
rect 10652 5176 10658 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11241 5219 11299 5225
rect 11241 5185 11253 5219
rect 11287 5216 11299 5219
rect 11514 5216 11520 5228
rect 11287 5188 11520 5216
rect 11287 5185 11299 5188
rect 11241 5179 11299 5185
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 12544 5225 12572 5256
rect 12636 5228 12664 5324
rect 12710 5312 12716 5364
rect 12768 5312 12774 5364
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 13722 5352 13728 5364
rect 13504 5324 13728 5352
rect 13504 5312 13510 5324
rect 13722 5312 13728 5324
rect 13780 5352 13786 5364
rect 15289 5355 15347 5361
rect 13780 5324 14228 5352
rect 13780 5312 13786 5324
rect 12728 5284 12756 5312
rect 13817 5287 13875 5293
rect 12728 5256 13584 5284
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 9858 5108 9864 5160
rect 9916 5108 9922 5160
rect 10686 5108 10692 5160
rect 10744 5108 10750 5160
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5117 10931 5151
rect 10873 5111 10931 5117
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 9950 5040 9956 5092
rect 10008 5080 10014 5092
rect 10781 5083 10839 5089
rect 10781 5080 10793 5083
rect 10008 5052 10793 5080
rect 10008 5040 10014 5052
rect 10781 5049 10793 5052
rect 10827 5049 10839 5083
rect 10888 5080 10916 5111
rect 11422 5080 11428 5092
rect 10888 5052 11428 5080
rect 10781 5043 10839 5049
rect 11422 5040 11428 5052
rect 11480 5040 11486 5092
rect 11992 5080 12020 5111
rect 12066 5108 12072 5160
rect 12124 5108 12130 5160
rect 12544 5080 12572 5179
rect 12618 5176 12624 5228
rect 12676 5176 12682 5228
rect 12802 5176 12808 5228
rect 12860 5176 12866 5228
rect 12894 5176 12900 5228
rect 12952 5216 12958 5228
rect 13556 5225 13584 5256
rect 13817 5253 13829 5287
rect 13863 5284 13875 5287
rect 14090 5284 14096 5296
rect 13863 5256 14096 5284
rect 13863 5253 13875 5256
rect 13817 5247 13875 5253
rect 14090 5244 14096 5256
rect 14148 5244 14154 5296
rect 14200 5284 14228 5324
rect 15289 5321 15301 5355
rect 15335 5352 15347 5355
rect 15378 5352 15384 5364
rect 15335 5324 15384 5352
rect 15335 5321 15347 5324
rect 15289 5315 15347 5321
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 14200 5256 14306 5284
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12952 5188 13001 5216
rect 12952 5176 12958 5188
rect 12989 5185 13001 5188
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5148 12771 5151
rect 12912 5148 12940 5176
rect 13096 5148 13124 5179
rect 12759 5120 12940 5148
rect 13004 5120 13124 5148
rect 12759 5117 12771 5120
rect 12713 5111 12771 5117
rect 13004 5080 13032 5120
rect 11992 5052 12112 5080
rect 12544 5052 13032 5080
rect 12084 5024 12112 5052
rect 10962 5012 10968 5024
rect 9646 4984 10968 5012
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11146 4972 11152 5024
rect 11204 4972 11210 5024
rect 12066 4972 12072 5024
rect 12124 5012 12130 5024
rect 12345 5015 12403 5021
rect 12345 5012 12357 5015
rect 12124 4984 12357 5012
rect 12124 4972 12130 4984
rect 12345 4981 12357 4984
rect 12391 4981 12403 5015
rect 12345 4975 12403 4981
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12805 5015 12863 5021
rect 12805 5012 12817 5015
rect 12584 4984 12817 5012
rect 12584 4972 12590 4984
rect 12805 4981 12817 4984
rect 12851 4981 12863 5015
rect 12805 4975 12863 4981
rect 1104 4922 16008 4944
rect 1104 4870 2813 4922
rect 2865 4870 2877 4922
rect 2929 4870 2941 4922
rect 2993 4870 3005 4922
rect 3057 4870 3069 4922
rect 3121 4870 6539 4922
rect 6591 4870 6603 4922
rect 6655 4870 6667 4922
rect 6719 4870 6731 4922
rect 6783 4870 6795 4922
rect 6847 4870 10265 4922
rect 10317 4870 10329 4922
rect 10381 4870 10393 4922
rect 10445 4870 10457 4922
rect 10509 4870 10521 4922
rect 10573 4870 13991 4922
rect 14043 4870 14055 4922
rect 14107 4870 14119 4922
rect 14171 4870 14183 4922
rect 14235 4870 14247 4922
rect 14299 4870 16008 4922
rect 1104 4848 16008 4870
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3786 4808 3792 4820
rect 3651 4780 3792 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4065 4811 4123 4817
rect 4065 4777 4077 4811
rect 4111 4808 4123 4811
rect 4338 4808 4344 4820
rect 4111 4780 4344 4808
rect 4111 4777 4123 4780
rect 4065 4771 4123 4777
rect 4338 4768 4344 4780
rect 4396 4768 4402 4820
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 4801 4811 4859 4817
rect 4801 4808 4813 4811
rect 4672 4780 4813 4808
rect 4672 4768 4678 4780
rect 4801 4777 4813 4780
rect 4847 4777 4859 4811
rect 4801 4771 4859 4777
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 4985 4811 5043 4817
rect 4985 4808 4997 4811
rect 4948 4780 4997 4808
rect 4948 4768 4954 4780
rect 4985 4777 4997 4780
rect 5031 4777 5043 4811
rect 4985 4771 5043 4777
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5224 4780 5273 4808
rect 5224 4768 5230 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 5353 4811 5411 4817
rect 5353 4777 5365 4811
rect 5399 4808 5411 4811
rect 5994 4808 6000 4820
rect 5399 4780 6000 4808
rect 5399 4777 5411 4780
rect 5353 4771 5411 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6086 4768 6092 4820
rect 6144 4768 6150 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7248 4780 8708 4808
rect 7248 4768 7254 4780
rect 4430 4740 4436 4752
rect 4080 4712 4436 4740
rect 1854 4632 1860 4684
rect 1912 4632 1918 4684
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4672 2191 4675
rect 2498 4672 2504 4684
rect 2179 4644 2504 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3418 4604 3424 4616
rect 3292 4576 3424 4604
rect 3292 4564 3298 4576
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 4080 4613 4108 4712
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 4632 4672 4660 4768
rect 4264 4644 4660 4672
rect 4264 4613 4292 4644
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 5169 4675 5227 4681
rect 5169 4672 5181 4675
rect 4764 4644 5181 4672
rect 4764 4632 4770 4644
rect 5169 4641 5181 4644
rect 5215 4641 5227 4675
rect 6104 4672 6132 4768
rect 8389 4743 8447 4749
rect 8389 4709 8401 4743
rect 8435 4709 8447 4743
rect 8389 4703 8447 4709
rect 5169 4635 5227 4641
rect 5460 4644 6132 4672
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 3804 4536 3832 4567
rect 4356 4536 4384 4567
rect 3804 4508 4384 4536
rect 4080 4480 4108 4508
rect 4062 4428 4068 4480
rect 4120 4428 4126 4480
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4540 4468 4568 4567
rect 4614 4564 4620 4616
rect 4672 4604 4678 4616
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 4672 4576 4905 4604
rect 4672 4564 4678 4576
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 4982 4564 4988 4616
rect 5040 4604 5046 4616
rect 5460 4613 5488 4644
rect 6270 4632 6276 4684
rect 6328 4672 6334 4684
rect 6549 4675 6607 4681
rect 6549 4672 6561 4675
rect 6328 4644 6561 4672
rect 6328 4632 6334 4644
rect 6549 4641 6561 4644
rect 6595 4641 6607 4675
rect 6549 4635 6607 4641
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 8404 4672 8432 4703
rect 6871 4644 8432 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 5077 4607 5135 4613
rect 5077 4604 5089 4607
rect 5040 4576 5089 4604
rect 5040 4564 5046 4576
rect 5077 4573 5089 4576
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 6086 4564 6092 4616
rect 6144 4564 6150 4616
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 7892 4576 7958 4604
rect 7892 4564 7898 4576
rect 8294 4564 8300 4616
rect 8352 4604 8358 4616
rect 8680 4613 8708 4780
rect 10686 4768 10692 4820
rect 10744 4768 10750 4820
rect 12529 4811 12587 4817
rect 12529 4808 12541 4811
rect 11256 4780 12541 4808
rect 11256 4740 11284 4780
rect 12529 4777 12541 4780
rect 12575 4808 12587 4811
rect 12802 4808 12808 4820
rect 12575 4780 12808 4808
rect 12575 4777 12587 4780
rect 12529 4771 12587 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 13906 4768 13912 4820
rect 13964 4808 13970 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13964 4780 14105 4808
rect 13964 4768 13970 4780
rect 14093 4777 14105 4780
rect 14139 4808 14151 4811
rect 14274 4808 14280 4820
rect 14139 4780 14280 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 14829 4811 14887 4817
rect 14829 4808 14841 4811
rect 14424 4780 14841 4808
rect 14424 4768 14430 4780
rect 10796 4712 11284 4740
rect 8938 4632 8944 4684
rect 8996 4632 9002 4684
rect 9214 4632 9220 4684
rect 9272 4632 9278 4684
rect 10796 4616 10824 4712
rect 11514 4700 11520 4752
rect 11572 4740 11578 4752
rect 13633 4743 13691 4749
rect 11572 4712 12572 4740
rect 11572 4700 11578 4712
rect 10962 4632 10968 4684
rect 11020 4632 11026 4684
rect 11440 4644 12388 4672
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 8352 4576 8401 4604
rect 8352 4564 8358 4576
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4573 8723 4607
rect 8665 4567 8723 4573
rect 10778 4564 10784 4616
rect 10836 4564 10842 4616
rect 11146 4564 11152 4616
rect 11204 4604 11210 4616
rect 11204 4600 11284 4604
rect 11440 4600 11468 4644
rect 11204 4576 11468 4600
rect 11204 4564 11210 4576
rect 11256 4572 11468 4576
rect 11514 4564 11520 4616
rect 11572 4564 11578 4616
rect 12360 4613 12388 4644
rect 12544 4613 12572 4712
rect 13633 4709 13645 4743
rect 13679 4709 13691 4743
rect 13633 4703 13691 4709
rect 13081 4675 13139 4681
rect 13081 4641 13093 4675
rect 13127 4672 13139 4675
rect 13127 4644 13584 4672
rect 13127 4641 13139 4644
rect 13081 4635 13139 4641
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 10502 4536 10508 4548
rect 4632 4508 7236 4536
rect 4632 4477 4660 4508
rect 4212 4440 4568 4468
rect 4617 4471 4675 4477
rect 4212 4428 4218 4440
rect 4617 4437 4629 4471
rect 4663 4437 4675 4471
rect 4617 4431 4675 4437
rect 5534 4428 5540 4480
rect 5592 4428 5598 4480
rect 7208 4468 7236 4508
rect 8220 4508 9628 4536
rect 10442 4508 10508 4536
rect 8220 4468 8248 4508
rect 7208 4440 8248 4468
rect 8294 4428 8300 4480
rect 8352 4428 8358 4480
rect 8570 4428 8576 4480
rect 8628 4428 8634 4480
rect 9600 4468 9628 4508
rect 10502 4496 10508 4508
rect 10560 4536 10566 4548
rect 10686 4536 10692 4548
rect 10560 4508 10692 4536
rect 10560 4496 10566 4508
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 12176 4536 12204 4567
rect 11440 4508 12204 4536
rect 12360 4536 12388 4567
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 13265 4607 13323 4613
rect 13265 4604 13277 4607
rect 12676 4576 13277 4604
rect 12676 4564 12682 4576
rect 13265 4573 13277 4576
rect 13311 4573 13323 4607
rect 13265 4567 13323 4573
rect 13556 4536 13584 4644
rect 13648 4604 13676 4703
rect 13909 4607 13967 4613
rect 13909 4604 13921 4607
rect 13648 4576 13921 4604
rect 13909 4573 13921 4576
rect 13955 4573 13967 4607
rect 13909 4567 13967 4573
rect 13998 4564 14004 4616
rect 14056 4604 14062 4616
rect 14476 4613 14504 4780
rect 14829 4777 14841 4780
rect 14875 4777 14887 4811
rect 14829 4771 14887 4777
rect 14645 4675 14703 4681
rect 14645 4641 14657 4675
rect 14691 4672 14703 4675
rect 14691 4644 15148 4672
rect 14691 4641 14703 4644
rect 14645 4635 14703 4641
rect 14277 4607 14335 4613
rect 14277 4604 14289 4607
rect 14056 4576 14289 4604
rect 14056 4564 14062 4576
rect 14277 4573 14289 4576
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 14090 4536 14096 4548
rect 12360 4508 13216 4536
rect 13556 4508 14096 4536
rect 11440 4480 11468 4508
rect 13188 4480 13216 4508
rect 14090 4496 14096 4508
rect 14148 4496 14154 4548
rect 14384 4536 14412 4567
rect 14660 4536 14688 4635
rect 15120 4616 15148 4644
rect 14921 4607 14979 4613
rect 14921 4573 14933 4607
rect 14967 4573 14979 4607
rect 14921 4567 14979 4573
rect 14384 4508 14688 4536
rect 14936 4536 14964 4567
rect 15010 4564 15016 4616
rect 15068 4564 15074 4616
rect 15102 4564 15108 4616
rect 15160 4564 15166 4616
rect 15470 4536 15476 4548
rect 14936 4508 15476 4536
rect 15470 4496 15476 4508
rect 15528 4496 15534 4548
rect 11330 4468 11336 4480
rect 9600 4440 11336 4468
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 11422 4428 11428 4480
rect 11480 4428 11486 4480
rect 11606 4428 11612 4480
rect 11664 4428 11670 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 12710 4468 12716 4480
rect 12492 4440 12716 4468
rect 12492 4428 12498 4440
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 13170 4428 13176 4480
rect 13228 4428 13234 4480
rect 13722 4428 13728 4480
rect 13780 4428 13786 4480
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 14240 4440 14657 4468
rect 14240 4428 14246 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 14645 4431 14703 4437
rect 15654 4428 15660 4480
rect 15712 4428 15718 4480
rect 1104 4378 16008 4400
rect 1104 4326 3473 4378
rect 3525 4326 3537 4378
rect 3589 4326 3601 4378
rect 3653 4326 3665 4378
rect 3717 4326 3729 4378
rect 3781 4326 7199 4378
rect 7251 4326 7263 4378
rect 7315 4326 7327 4378
rect 7379 4326 7391 4378
rect 7443 4326 7455 4378
rect 7507 4326 10925 4378
rect 10977 4326 10989 4378
rect 11041 4326 11053 4378
rect 11105 4326 11117 4378
rect 11169 4326 11181 4378
rect 11233 4326 14651 4378
rect 14703 4326 14715 4378
rect 14767 4326 14779 4378
rect 14831 4326 14843 4378
rect 14895 4326 14907 4378
rect 14959 4326 16008 4378
rect 1104 4304 16008 4326
rect 3605 4267 3663 4273
rect 3605 4233 3617 4267
rect 3651 4264 3663 4267
rect 3878 4264 3884 4276
rect 3651 4236 3884 4264
rect 3651 4233 3663 4236
rect 3605 4227 3663 4233
rect 3878 4224 3884 4236
rect 3936 4224 3942 4276
rect 4062 4224 4068 4276
rect 4120 4224 4126 4276
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 5442 4264 5448 4276
rect 4488 4236 5448 4264
rect 4488 4224 4494 4236
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 5997 4267 6055 4273
rect 5997 4233 6009 4267
rect 6043 4264 6055 4267
rect 6086 4264 6092 4276
rect 6043 4236 6092 4264
rect 6043 4233 6055 4236
rect 5997 4227 6055 4233
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 6932 4236 7788 4264
rect 3786 4196 3792 4208
rect 3712 4168 3792 4196
rect 1854 4088 1860 4140
rect 1912 4088 1918 4140
rect 3234 4088 3240 4140
rect 3292 4088 3298 4140
rect 3712 4137 3740 4168
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 3896 4196 3924 4224
rect 4614 4196 4620 4208
rect 3896 4168 4620 4196
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4128 3939 4131
rect 4062 4128 4068 4140
rect 3927 4100 4068 4128
rect 3927 4097 3939 4100
rect 3881 4091 3939 4097
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 3142 4060 3148 4072
rect 2179 4032 3148 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3326 4020 3332 4072
rect 3384 4060 3390 4072
rect 3789 4063 3847 4069
rect 3789 4060 3801 4063
rect 3384 4032 3801 4060
rect 3384 4020 3390 4032
rect 3789 4029 3801 4032
rect 3835 4029 3847 4063
rect 3789 4023 3847 4029
rect 3896 3992 3924 4091
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4172 4137 4200 4168
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 6932 4196 6960 4236
rect 5750 4168 6960 4196
rect 7760 4140 7788 4236
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 11241 4267 11299 4273
rect 9180 4236 11100 4264
rect 9180 4224 9186 4236
rect 11072 4196 11100 4236
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11422 4264 11428 4276
rect 11287 4236 11428 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11422 4224 11428 4236
rect 11480 4224 11486 4276
rect 14182 4264 14188 4276
rect 12452 4236 14188 4264
rect 11885 4199 11943 4205
rect 11885 4196 11897 4199
rect 11072 4168 11897 4196
rect 11885 4165 11897 4168
rect 11931 4165 11943 4199
rect 11885 4159 11943 4165
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 6270 4088 6276 4140
rect 6328 4128 6334 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 6328 4100 6377 4128
rect 6328 4088 6334 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 8352 4100 8493 4128
rect 8352 4088 8358 4100
rect 8481 4097 8493 4100
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9490 4128 9496 4140
rect 8996 4100 9496 4128
rect 8996 4088 9002 4100
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 10902 4114 11100 4128
rect 10888 4100 11100 4114
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 3344 3964 3924 3992
rect 3344 3936 3372 3964
rect 3326 3884 3332 3936
rect 3384 3884 3390 3936
rect 4264 3924 4292 4023
rect 4522 4020 4528 4072
rect 4580 4020 4586 4072
rect 6288 3992 6316 4088
rect 6641 4063 6699 4069
rect 6641 4060 6653 4063
rect 5552 3964 6316 3992
rect 6380 4032 6653 4060
rect 5552 3924 5580 3964
rect 4264 3896 5580 3924
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6380 3924 6408 4032
rect 6641 4029 6653 4032
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8628 4032 9137 4060
rect 8628 4020 8634 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9766 4020 9772 4072
rect 9824 4020 9830 4072
rect 10502 4020 10508 4072
rect 10560 4060 10566 4072
rect 10888 4060 10916 4100
rect 10560 4032 10916 4060
rect 11072 4060 11100 4100
rect 11330 4088 11336 4140
rect 11388 4128 11394 4140
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 11388 4100 11805 4128
rect 11388 4088 11394 4100
rect 11793 4097 11805 4100
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12452 4128 12480 4236
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 14274 4224 14280 4276
rect 14332 4264 14338 4276
rect 14737 4267 14795 4273
rect 14737 4264 14749 4267
rect 14332 4236 14749 4264
rect 14332 4224 14338 4236
rect 14737 4233 14749 4236
rect 14783 4264 14795 4267
rect 15010 4264 15016 4276
rect 14783 4236 15016 4264
rect 14783 4233 14795 4236
rect 14737 4227 14795 4233
rect 15010 4224 15016 4236
rect 15068 4224 15074 4276
rect 15470 4224 15476 4276
rect 15528 4224 15534 4276
rect 12710 4196 12716 4208
rect 12544 4168 12716 4196
rect 12544 4137 12572 4168
rect 12710 4156 12716 4168
rect 12768 4156 12774 4208
rect 13906 4156 13912 4208
rect 13964 4156 13970 4208
rect 12023 4100 12480 4128
rect 12529 4131 12587 4137
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 11072 4032 11376 4060
rect 10560 4020 10566 4032
rect 11348 4004 11376 4032
rect 11514 4020 11520 4072
rect 11572 4020 11578 4072
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 12345 4063 12403 4069
rect 12345 4060 12357 4063
rect 11756 4032 12357 4060
rect 11756 4020 11762 4032
rect 12345 4029 12357 4032
rect 12391 4029 12403 4063
rect 12345 4023 12403 4029
rect 12434 4020 12440 4072
rect 12492 4060 12498 4072
rect 12544 4060 12572 4091
rect 12618 4088 12624 4140
rect 12676 4088 12682 4140
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12860 4100 12909 4128
rect 12860 4088 12866 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 14550 4088 14556 4140
rect 14608 4128 14614 4140
rect 15013 4131 15071 4137
rect 15013 4128 15025 4131
rect 14608 4100 15025 4128
rect 14608 4088 14614 4100
rect 15013 4097 15025 4100
rect 15059 4097 15071 4131
rect 15381 4131 15439 4137
rect 15381 4128 15393 4131
rect 15013 4091 15071 4097
rect 15120 4100 15393 4128
rect 12492 4032 12572 4060
rect 13265 4063 13323 4069
rect 12492 4020 12498 4032
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13722 4060 13728 4072
rect 13311 4032 13728 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14458 4020 14464 4072
rect 14516 4060 14522 4072
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 14516 4032 14841 4060
rect 14516 4020 14522 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 14918 4020 14924 4072
rect 14976 4060 14982 4072
rect 15120 4060 15148 4100
rect 15381 4097 15393 4100
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 14976 4032 15148 4060
rect 14976 4020 14982 4032
rect 15286 4020 15292 4072
rect 15344 4020 15350 4072
rect 11330 3952 11336 4004
rect 11388 3952 11394 4004
rect 11609 3995 11667 4001
rect 11609 3961 11621 3995
rect 11655 3992 11667 3995
rect 12158 3992 12164 4004
rect 11655 3964 12164 3992
rect 11655 3961 11667 3964
rect 11609 3955 11667 3961
rect 12158 3952 12164 3964
rect 12216 3952 12222 4004
rect 12253 3995 12311 4001
rect 12253 3961 12265 3995
rect 12299 3992 12311 3995
rect 12710 3992 12716 4004
rect 12299 3964 12716 3992
rect 12299 3961 12311 3964
rect 12253 3955 12311 3961
rect 12710 3952 12716 3964
rect 12768 3952 12774 4004
rect 15197 3995 15255 4001
rect 15197 3992 15209 3995
rect 14292 3964 15209 3992
rect 6144 3896 6408 3924
rect 6144 3884 6150 3896
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 8113 3927 8171 3933
rect 8113 3924 8125 3927
rect 6512 3896 8125 3924
rect 6512 3884 6518 3896
rect 8113 3893 8125 3896
rect 8159 3893 8171 3927
rect 8113 3887 8171 3893
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 12805 3927 12863 3933
rect 12805 3924 12817 3927
rect 8352 3896 12817 3924
rect 8352 3884 8358 3896
rect 12805 3893 12817 3896
rect 12851 3924 12863 3927
rect 14292 3924 14320 3964
rect 15197 3961 15209 3964
rect 15243 3961 15255 3995
rect 15197 3955 15255 3961
rect 12851 3896 14320 3924
rect 12851 3893 12863 3896
rect 12805 3887 12863 3893
rect 1104 3834 16008 3856
rect 1104 3782 2813 3834
rect 2865 3782 2877 3834
rect 2929 3782 2941 3834
rect 2993 3782 3005 3834
rect 3057 3782 3069 3834
rect 3121 3782 6539 3834
rect 6591 3782 6603 3834
rect 6655 3782 6667 3834
rect 6719 3782 6731 3834
rect 6783 3782 6795 3834
rect 6847 3782 10265 3834
rect 10317 3782 10329 3834
rect 10381 3782 10393 3834
rect 10445 3782 10457 3834
rect 10509 3782 10521 3834
rect 10573 3782 13991 3834
rect 14043 3782 14055 3834
rect 14107 3782 14119 3834
rect 14171 3782 14183 3834
rect 14235 3782 14247 3834
rect 14299 3782 16008 3834
rect 1104 3760 16008 3782
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 4893 3723 4951 3729
rect 4893 3720 4905 3723
rect 4580 3692 4905 3720
rect 4580 3680 4586 3692
rect 4893 3689 4905 3692
rect 4939 3689 4951 3723
rect 4893 3683 4951 3689
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5721 3723 5779 3729
rect 5721 3720 5733 3723
rect 5592 3692 5733 3720
rect 5592 3680 5598 3692
rect 5721 3689 5733 3692
rect 5767 3689 5779 3723
rect 5721 3683 5779 3689
rect 6086 3680 6092 3732
rect 6144 3680 6150 3732
rect 6270 3680 6276 3732
rect 6328 3680 6334 3732
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 7926 3720 7932 3732
rect 7708 3692 7932 3720
rect 7708 3680 7714 3692
rect 7926 3680 7932 3692
rect 7984 3680 7990 3732
rect 9309 3723 9367 3729
rect 9309 3689 9321 3723
rect 9355 3720 9367 3723
rect 9858 3720 9864 3732
rect 9355 3692 9864 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 9950 3680 9956 3732
rect 10008 3680 10014 3732
rect 10216 3723 10274 3729
rect 10216 3689 10228 3723
rect 10262 3720 10274 3723
rect 11698 3720 11704 3732
rect 10262 3692 11704 3720
rect 10262 3689 10274 3692
rect 10216 3683 10274 3689
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 13630 3680 13636 3732
rect 13688 3680 13694 3732
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 14918 3720 14924 3732
rect 13964 3692 14924 3720
rect 13964 3680 13970 3692
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 15286 3680 15292 3732
rect 15344 3680 15350 3732
rect 4982 3652 4988 3664
rect 4356 3624 4988 3652
rect 1854 3544 1860 3596
rect 1912 3544 1918 3596
rect 4356 3593 4384 3624
rect 4982 3612 4988 3624
rect 5040 3612 5046 3664
rect 3605 3587 3663 3593
rect 3605 3553 3617 3587
rect 3651 3584 3663 3587
rect 4341 3587 4399 3593
rect 4341 3584 4353 3587
rect 3651 3556 4353 3584
rect 3651 3553 3663 3556
rect 3605 3547 3663 3553
rect 4341 3553 4353 3556
rect 4387 3553 4399 3587
rect 4341 3547 4399 3553
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3584 4859 3587
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 4847 3556 5273 3584
rect 4847 3553 4859 3556
rect 4801 3547 4859 3553
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5261 3547 5319 3553
rect 3234 3476 3240 3528
rect 3292 3476 3298 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3516 5135 3519
rect 5169 3519 5227 3525
rect 5169 3516 5181 3519
rect 5123 3488 5181 3516
rect 5123 3485 5135 3488
rect 5077 3479 5135 3485
rect 5169 3485 5181 3488
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5442 3516 5448 3528
rect 5399 3488 5448 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 2130 3408 2136 3460
rect 2188 3408 2194 3460
rect 3789 3383 3847 3389
rect 3789 3349 3801 3383
rect 3835 3380 3847 3383
rect 3878 3380 3884 3392
rect 3835 3352 3884 3380
rect 3835 3349 3847 3352
rect 3789 3343 3847 3349
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 5000 3380 5028 3479
rect 5184 3448 5212 3479
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 5552 3448 5580 3680
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3584 6239 3587
rect 6288 3584 6316 3680
rect 9968 3652 9996 3680
rect 9416 3624 9996 3652
rect 9416 3593 9444 3624
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 11885 3655 11943 3661
rect 11885 3652 11897 3655
rect 11572 3624 11897 3652
rect 11572 3612 11578 3624
rect 11885 3621 11897 3624
rect 11931 3621 11943 3655
rect 11885 3615 11943 3621
rect 6227 3556 6316 3584
rect 6457 3587 6515 3593
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 6457 3553 6469 3587
rect 6503 3584 6515 3587
rect 8665 3587 8723 3593
rect 8665 3584 8677 3587
rect 6503 3556 8677 3584
rect 6503 3553 6515 3556
rect 6457 3547 6515 3553
rect 8665 3553 8677 3556
rect 8711 3553 8723 3587
rect 9401 3587 9459 3593
rect 8665 3547 8723 3553
rect 9140 3556 9352 3584
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 5902 3476 5908 3528
rect 5960 3476 5966 3528
rect 7742 3516 7748 3528
rect 7590 3488 7748 3516
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7984 3488 8217 3516
rect 7984 3476 7990 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8294 3476 8300 3528
rect 8352 3476 8358 3528
rect 9140 3525 9168 3556
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3485 9275 3519
rect 9324 3516 9352 3556
rect 9401 3553 9413 3587
rect 9447 3553 9459 3587
rect 9401 3547 9459 3553
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9548 3556 9965 3584
rect 9548 3544 9554 3556
rect 9953 3553 9965 3556
rect 9999 3584 10011 3587
rect 12161 3587 12219 3593
rect 12161 3584 12173 3587
rect 9999 3556 12173 3584
rect 9999 3553 10011 3556
rect 9953 3547 10011 3553
rect 12161 3553 12173 3556
rect 12207 3584 12219 3587
rect 12986 3584 12992 3596
rect 12207 3556 12992 3584
rect 12207 3553 12219 3556
rect 12161 3547 12219 3553
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 9324 3488 9996 3516
rect 9217 3479 9275 3485
rect 5184 3420 5580 3448
rect 5166 3380 5172 3392
rect 5000 3352 5172 3380
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 5920 3380 5948 3476
rect 8496 3448 8524 3479
rect 9232 3448 9260 3479
rect 7852 3420 9260 3448
rect 9968 3448 9996 3488
rect 11330 3476 11336 3528
rect 11388 3476 11394 3528
rect 11974 3516 11980 3528
rect 11716 3488 11980 3516
rect 9968 3420 10640 3448
rect 7852 3380 7880 3420
rect 10612 3392 10640 3420
rect 5920 3352 7880 3380
rect 10594 3340 10600 3392
rect 10652 3340 10658 3392
rect 11716 3389 11744 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 13648 3516 13676 3680
rect 15304 3652 15332 3680
rect 15473 3655 15531 3661
rect 15473 3652 15485 3655
rect 15304 3624 15485 3652
rect 15473 3621 15485 3624
rect 15519 3621 15531 3655
rect 15473 3615 15531 3621
rect 13998 3516 14004 3528
rect 13570 3488 14004 3516
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 14921 3519 14979 3525
rect 14921 3485 14933 3519
rect 14967 3516 14979 3519
rect 15102 3516 15108 3528
rect 14967 3488 15108 3516
rect 14967 3485 14979 3488
rect 14921 3479 14979 3485
rect 12437 3451 12495 3457
rect 12437 3417 12449 3451
rect 12483 3417 12495 3451
rect 14093 3451 14151 3457
rect 14093 3448 14105 3451
rect 12437 3411 12495 3417
rect 13740 3420 14105 3448
rect 11701 3383 11759 3389
rect 11701 3349 11713 3383
rect 11747 3349 11759 3383
rect 12452 3380 12480 3411
rect 13740 3380 13768 3420
rect 14093 3417 14105 3420
rect 14139 3417 14151 3451
rect 14752 3448 14780 3479
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 15010 3448 15016 3460
rect 14752 3420 15016 3448
rect 14093 3411 14151 3417
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 12452 3352 13768 3380
rect 11701 3343 11759 3349
rect 1104 3290 16008 3312
rect 1104 3238 3473 3290
rect 3525 3238 3537 3290
rect 3589 3238 3601 3290
rect 3653 3238 3665 3290
rect 3717 3238 3729 3290
rect 3781 3238 7199 3290
rect 7251 3238 7263 3290
rect 7315 3238 7327 3290
rect 7379 3238 7391 3290
rect 7443 3238 7455 3290
rect 7507 3238 10925 3290
rect 10977 3238 10989 3290
rect 11041 3238 11053 3290
rect 11105 3238 11117 3290
rect 11169 3238 11181 3290
rect 11233 3238 14651 3290
rect 14703 3238 14715 3290
rect 14767 3238 14779 3290
rect 14831 3238 14843 3290
rect 14895 3238 14907 3290
rect 14959 3238 16008 3290
rect 1104 3216 16008 3238
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 2869 3179 2927 3185
rect 2869 3176 2881 3179
rect 2188 3148 2881 3176
rect 2188 3136 2194 3148
rect 2869 3145 2881 3148
rect 2915 3145 2927 3179
rect 2869 3139 2927 3145
rect 3878 3136 3884 3188
rect 3936 3136 3942 3188
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 6457 3179 6515 3185
rect 6457 3176 6469 3179
rect 5684 3148 6469 3176
rect 5684 3136 5690 3148
rect 6457 3145 6469 3148
rect 6503 3145 6515 3179
rect 6457 3139 6515 3145
rect 7926 3136 7932 3188
rect 7984 3136 7990 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10229 3179 10287 3185
rect 10229 3176 10241 3179
rect 9824 3148 10241 3176
rect 9824 3136 9830 3148
rect 10229 3145 10241 3148
rect 10275 3145 10287 3179
rect 10229 3139 10287 3145
rect 10778 3136 10784 3188
rect 10836 3176 10842 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 10836 3148 10977 3176
rect 10836 3136 10842 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 10965 3139 11023 3145
rect 11974 3136 11980 3188
rect 12032 3136 12038 3188
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 12618 3176 12624 3188
rect 12124 3148 12624 3176
rect 12124 3136 12130 3148
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 12989 3179 13047 3185
rect 12989 3176 13001 3179
rect 12860 3148 13001 3176
rect 12860 3136 12866 3148
rect 12989 3145 13001 3148
rect 13035 3145 13047 3179
rect 14366 3176 14372 3188
rect 12989 3139 13047 3145
rect 13372 3148 14372 3176
rect 3326 3108 3332 3120
rect 3252 3080 3332 3108
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 3252 3049 3280 3080
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2832 3012 3065 3040
rect 2832 3000 2838 3012
rect 3053 3009 3065 3012
rect 3099 3009 3111 3043
rect 3053 3003 3111 3009
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3040 3571 3043
rect 3896 3040 3924 3136
rect 5902 3068 5908 3120
rect 5960 3108 5966 3120
rect 7944 3108 7972 3136
rect 5960 3080 7328 3108
rect 5960 3068 5966 3080
rect 3559 3012 3924 3040
rect 3559 3009 3571 3012
rect 3513 3003 3571 3009
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6512 3012 7021 3040
rect 6512 3000 6518 3012
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 1670 2932 1676 2984
rect 1728 2972 1734 2984
rect 3329 2975 3387 2981
rect 3329 2972 3341 2975
rect 1728 2944 3341 2972
rect 1728 2932 1734 2944
rect 3329 2941 3341 2944
rect 3375 2972 3387 2975
rect 7024 2972 7052 3003
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7300 3049 7328 3080
rect 7852 3080 7972 3108
rect 10428 3080 10732 3108
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 7156 3012 7205 3040
rect 7156 3000 7162 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 7285 3043 7343 3049
rect 7285 3009 7297 3043
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 7852 3049 7880 3080
rect 10428 3049 10456 3080
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 10413 3043 10471 3049
rect 10413 3009 10425 3043
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3009 10563 3043
rect 10505 3003 10563 3009
rect 7944 2972 7972 3003
rect 3375 2944 6960 2972
rect 7024 2944 7972 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 3145 2907 3203 2913
rect 3145 2873 3157 2907
rect 3191 2873 3203 2907
rect 6932 2904 6960 2944
rect 8294 2904 8300 2916
rect 6932 2876 8300 2904
rect 3145 2867 3203 2873
rect 3160 2836 3188 2867
rect 8294 2864 8300 2876
rect 8352 2864 8358 2916
rect 4430 2836 4436 2848
rect 3160 2808 4436 2836
rect 4430 2796 4436 2808
rect 4488 2796 4494 2848
rect 10520 2836 10548 3003
rect 10704 2972 10732 3080
rect 10796 3080 11652 3108
rect 10796 3049 10824 3080
rect 11624 3052 11652 3080
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3009 10839 3043
rect 10781 3003 10839 3009
rect 11057 3043 11115 3049
rect 11057 3009 11069 3043
rect 11103 3040 11115 3043
rect 11422 3040 11428 3052
rect 11103 3012 11428 3040
rect 11103 3009 11115 3012
rect 11057 3003 11115 3009
rect 11422 3000 11428 3012
rect 11480 3000 11486 3052
rect 11606 3000 11612 3052
rect 11664 3000 11670 3052
rect 11992 3040 12020 3136
rect 13372 3117 13400 3148
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 15010 3136 15016 3188
rect 15068 3136 15074 3188
rect 13357 3111 13415 3117
rect 13357 3077 13369 3111
rect 13403 3077 13415 3111
rect 13357 3071 13415 3077
rect 13998 3068 14004 3120
rect 14056 3068 14062 3120
rect 14921 3111 14979 3117
rect 14921 3077 14933 3111
rect 14967 3108 14979 3111
rect 15028 3108 15056 3136
rect 14967 3080 15056 3108
rect 14967 3077 14979 3080
rect 14921 3071 14979 3077
rect 12345 3043 12403 3049
rect 12345 3040 12357 3043
rect 11992 3012 12357 3040
rect 12345 3009 12357 3012
rect 12391 3009 12403 3043
rect 12345 3003 12403 3009
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 13081 3043 13139 3049
rect 13081 3040 13093 3043
rect 13044 3012 13093 3040
rect 13044 3000 13050 3012
rect 13081 3009 13093 3012
rect 13127 3009 13139 3043
rect 13081 3003 13139 3009
rect 15105 3043 15163 3049
rect 15105 3009 15117 3043
rect 15151 3009 15163 3043
rect 15105 3003 15163 3009
rect 15289 3043 15347 3049
rect 15289 3009 15301 3043
rect 15335 3040 15347 3043
rect 15654 3040 15660 3052
rect 15335 3012 15660 3040
rect 15335 3009 15347 3012
rect 15289 3003 15347 3009
rect 10704 2944 12434 2972
rect 10594 2864 10600 2916
rect 10652 2904 10658 2916
rect 10689 2907 10747 2913
rect 10689 2904 10701 2907
rect 10652 2876 10701 2904
rect 10652 2864 10658 2876
rect 10689 2873 10701 2876
rect 10735 2873 10747 2907
rect 10689 2867 10747 2873
rect 12406 2848 12434 2944
rect 13906 2932 13912 2984
rect 13964 2972 13970 2984
rect 13964 2944 14504 2972
rect 13964 2932 13970 2944
rect 14476 2904 14504 2944
rect 14550 2932 14556 2984
rect 14608 2972 14614 2984
rect 15120 2972 15148 3003
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 14608 2944 15148 2972
rect 15381 2975 15439 2981
rect 14608 2932 14614 2944
rect 15381 2941 15393 2975
rect 15427 2941 15439 2975
rect 15381 2935 15439 2941
rect 14734 2904 14740 2916
rect 14476 2876 14740 2904
rect 14734 2864 14740 2876
rect 14792 2904 14798 2916
rect 15396 2904 15424 2935
rect 14792 2876 15424 2904
rect 14792 2864 14798 2876
rect 12066 2836 12072 2848
rect 10520 2808 12072 2836
rect 12066 2796 12072 2808
rect 12124 2796 12130 2848
rect 12406 2808 12440 2848
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2836 14887 2839
rect 15102 2836 15108 2848
rect 14875 2808 15108 2836
rect 14875 2805 14887 2808
rect 14829 2799 14887 2805
rect 15102 2796 15108 2808
rect 15160 2796 15166 2848
rect 1104 2746 16008 2768
rect 1104 2694 2813 2746
rect 2865 2694 2877 2746
rect 2929 2694 2941 2746
rect 2993 2694 3005 2746
rect 3057 2694 3069 2746
rect 3121 2694 6539 2746
rect 6591 2694 6603 2746
rect 6655 2694 6667 2746
rect 6719 2694 6731 2746
rect 6783 2694 6795 2746
rect 6847 2694 10265 2746
rect 10317 2694 10329 2746
rect 10381 2694 10393 2746
rect 10445 2694 10457 2746
rect 10509 2694 10521 2746
rect 10573 2694 13991 2746
rect 14043 2694 14055 2746
rect 14107 2694 14119 2746
rect 14171 2694 14183 2746
rect 14235 2694 14247 2746
rect 14299 2694 16008 2746
rect 1104 2672 16008 2694
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 14645 2635 14703 2641
rect 14645 2632 14657 2635
rect 13228 2604 14657 2632
rect 13228 2592 13234 2604
rect 14645 2601 14657 2604
rect 14691 2601 14703 2635
rect 14645 2595 14703 2601
rect 1670 2524 1676 2576
rect 1728 2524 1734 2576
rect 14734 2524 14740 2576
rect 14792 2524 14798 2576
rect 15102 2456 15108 2508
rect 15160 2456 15166 2508
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 12710 2388 12716 2440
rect 12768 2428 12774 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12768 2400 13093 2428
rect 12768 2388 12774 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 72 2332 1501 2360
rect 72 2320 78 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1489 2323 1547 2329
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 9732 2264 9965 2292
rect 9732 2252 9738 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 9953 2255 10011 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 1104 2202 16008 2224
rect 1104 2150 3473 2202
rect 3525 2150 3537 2202
rect 3589 2150 3601 2202
rect 3653 2150 3665 2202
rect 3717 2150 3729 2202
rect 3781 2150 7199 2202
rect 7251 2150 7263 2202
rect 7315 2150 7327 2202
rect 7379 2150 7391 2202
rect 7443 2150 7455 2202
rect 7507 2150 10925 2202
rect 10977 2150 10989 2202
rect 11041 2150 11053 2202
rect 11105 2150 11117 2202
rect 11169 2150 11181 2202
rect 11233 2150 14651 2202
rect 14703 2150 14715 2202
rect 14767 2150 14779 2202
rect 14831 2150 14843 2202
rect 14895 2150 14907 2202
rect 14959 2150 16008 2202
rect 1104 2128 16008 2150
<< via1 >>
rect 2813 16838 2865 16890
rect 2877 16838 2929 16890
rect 2941 16838 2993 16890
rect 3005 16838 3057 16890
rect 3069 16838 3121 16890
rect 6539 16838 6591 16890
rect 6603 16838 6655 16890
rect 6667 16838 6719 16890
rect 6731 16838 6783 16890
rect 6795 16838 6847 16890
rect 10265 16838 10317 16890
rect 10329 16838 10381 16890
rect 10393 16838 10445 16890
rect 10457 16838 10509 16890
rect 10521 16838 10573 16890
rect 13991 16838 14043 16890
rect 14055 16838 14107 16890
rect 14119 16838 14171 16890
rect 14183 16838 14235 16890
rect 14247 16838 14299 16890
rect 8116 16600 8168 16652
rect 8392 16643 8444 16652
rect 8392 16609 8401 16643
rect 8401 16609 8435 16643
rect 8435 16609 8444 16643
rect 8392 16600 8444 16609
rect 11428 16600 11480 16652
rect 12900 16600 12952 16652
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 7656 16575 7708 16584
rect 7656 16541 7665 16575
rect 7665 16541 7699 16575
rect 7699 16541 7708 16575
rect 7656 16532 7708 16541
rect 11336 16532 11388 16584
rect 12348 16532 12400 16584
rect 4344 16396 4396 16448
rect 7104 16396 7156 16448
rect 9128 16396 9180 16448
rect 10784 16396 10836 16448
rect 3473 16294 3525 16346
rect 3537 16294 3589 16346
rect 3601 16294 3653 16346
rect 3665 16294 3717 16346
rect 3729 16294 3781 16346
rect 7199 16294 7251 16346
rect 7263 16294 7315 16346
rect 7327 16294 7379 16346
rect 7391 16294 7443 16346
rect 7455 16294 7507 16346
rect 10925 16294 10977 16346
rect 10989 16294 11041 16346
rect 11053 16294 11105 16346
rect 11117 16294 11169 16346
rect 11181 16294 11233 16346
rect 14651 16294 14703 16346
rect 14715 16294 14767 16346
rect 14779 16294 14831 16346
rect 14843 16294 14895 16346
rect 14907 16294 14959 16346
rect 4988 16235 5040 16244
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 5356 16192 5408 16244
rect 7104 16192 7156 16244
rect 9128 16192 9180 16244
rect 11428 16192 11480 16244
rect 6000 16056 6052 16108
rect 10140 16124 10192 16176
rect 10784 16124 10836 16176
rect 12440 16124 12492 16176
rect 12900 16099 12952 16108
rect 12900 16065 12909 16099
rect 12909 16065 12943 16099
rect 12943 16065 12952 16099
rect 12900 16056 12952 16065
rect 3884 15988 3936 16040
rect 5540 15988 5592 16040
rect 7932 16031 7984 16040
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 8208 16031 8260 16040
rect 8208 15997 8217 16031
rect 8217 15997 8251 16031
rect 8251 15997 8260 16031
rect 8208 15988 8260 15997
rect 12348 15988 12400 16040
rect 4620 15852 4672 15904
rect 5080 15895 5132 15904
rect 5080 15861 5089 15895
rect 5089 15861 5123 15895
rect 5123 15861 5132 15895
rect 5080 15852 5132 15861
rect 7840 15852 7892 15904
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 2813 15750 2865 15802
rect 2877 15750 2929 15802
rect 2941 15750 2993 15802
rect 3005 15750 3057 15802
rect 3069 15750 3121 15802
rect 6539 15750 6591 15802
rect 6603 15750 6655 15802
rect 6667 15750 6719 15802
rect 6731 15750 6783 15802
rect 6795 15750 6847 15802
rect 10265 15750 10317 15802
rect 10329 15750 10381 15802
rect 10393 15750 10445 15802
rect 10457 15750 10509 15802
rect 10521 15750 10573 15802
rect 13991 15750 14043 15802
rect 14055 15750 14107 15802
rect 14119 15750 14171 15802
rect 14183 15750 14235 15802
rect 14247 15750 14299 15802
rect 5080 15648 5132 15700
rect 7840 15648 7892 15700
rect 8208 15648 8260 15700
rect 10140 15648 10192 15700
rect 4620 15555 4672 15564
rect 4620 15521 4629 15555
rect 4629 15521 4663 15555
rect 4663 15521 4672 15555
rect 4620 15512 4672 15521
rect 7932 15512 7984 15564
rect 3148 15376 3200 15428
rect 2780 15308 2832 15360
rect 6000 15444 6052 15496
rect 6920 15444 6972 15496
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 9772 15444 9824 15496
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 11428 15512 11480 15564
rect 12164 15512 12216 15564
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 12900 15648 12952 15700
rect 4252 15308 4304 15360
rect 5632 15308 5684 15360
rect 6368 15351 6420 15360
rect 6368 15317 6377 15351
rect 6377 15317 6411 15351
rect 6411 15317 6420 15351
rect 6368 15308 6420 15317
rect 6552 15308 6604 15360
rect 9680 15351 9732 15360
rect 9680 15317 9689 15351
rect 9689 15317 9723 15351
rect 9723 15317 9732 15351
rect 9680 15308 9732 15317
rect 12900 15444 12952 15496
rect 11980 15308 12032 15360
rect 13268 15308 13320 15360
rect 13452 15351 13504 15360
rect 13452 15317 13461 15351
rect 13461 15317 13495 15351
rect 13495 15317 13504 15351
rect 13452 15308 13504 15317
rect 3473 15206 3525 15258
rect 3537 15206 3589 15258
rect 3601 15206 3653 15258
rect 3665 15206 3717 15258
rect 3729 15206 3781 15258
rect 7199 15206 7251 15258
rect 7263 15206 7315 15258
rect 7327 15206 7379 15258
rect 7391 15206 7443 15258
rect 7455 15206 7507 15258
rect 10925 15206 10977 15258
rect 10989 15206 11041 15258
rect 11053 15206 11105 15258
rect 11117 15206 11169 15258
rect 11181 15206 11233 15258
rect 14651 15206 14703 15258
rect 14715 15206 14767 15258
rect 14779 15206 14831 15258
rect 14843 15206 14895 15258
rect 14907 15206 14959 15258
rect 3884 15147 3936 15156
rect 3884 15113 3893 15147
rect 3893 15113 3927 15147
rect 3927 15113 3936 15147
rect 3884 15104 3936 15113
rect 3976 14968 4028 15020
rect 2780 14875 2832 14884
rect 2780 14841 2789 14875
rect 2789 14841 2823 14875
rect 2823 14841 2832 14875
rect 2780 14832 2832 14841
rect 2688 14764 2740 14816
rect 4252 15011 4304 15020
rect 4252 14977 4261 15011
rect 4261 14977 4295 15011
rect 4295 14977 4304 15011
rect 4252 14968 4304 14977
rect 4620 15036 4672 15088
rect 4988 15036 5040 15088
rect 6368 15104 6420 15156
rect 7656 15104 7708 15156
rect 7380 15036 7432 15088
rect 6000 14968 6052 15020
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 8392 15104 8444 15156
rect 8484 15104 8536 15156
rect 9128 15104 9180 15156
rect 6552 14968 6604 14977
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 4344 14943 4396 14952
rect 4344 14909 4353 14943
rect 4353 14909 4387 14943
rect 4387 14909 4396 14943
rect 4344 14900 4396 14909
rect 4712 14943 4764 14952
rect 4712 14909 4721 14943
rect 4721 14909 4755 14943
rect 4755 14909 4764 14943
rect 4712 14900 4764 14909
rect 5264 14764 5316 14816
rect 5448 14764 5500 14816
rect 7472 14900 7524 14952
rect 12900 15104 12952 15156
rect 9680 15079 9732 15088
rect 9680 15045 9689 15079
rect 9689 15045 9723 15079
rect 9723 15045 9732 15079
rect 9680 15036 9732 15045
rect 9772 15036 9824 15088
rect 10140 15036 10192 15088
rect 12716 15036 12768 15088
rect 14464 15104 14516 15156
rect 11980 14943 12032 14952
rect 6184 14807 6236 14816
rect 6184 14773 6193 14807
rect 6193 14773 6227 14807
rect 6227 14773 6236 14807
rect 6184 14764 6236 14773
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 9496 14764 9548 14816
rect 11980 14909 11989 14943
rect 11989 14909 12023 14943
rect 12023 14909 12032 14943
rect 11980 14900 12032 14909
rect 12256 14943 12308 14952
rect 12256 14909 12265 14943
rect 12265 14909 12299 14943
rect 12299 14909 12308 14943
rect 12256 14900 12308 14909
rect 15292 14943 15344 14952
rect 15292 14909 15301 14943
rect 15301 14909 15335 14943
rect 15335 14909 15344 14943
rect 15292 14900 15344 14909
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 11336 14764 11388 14816
rect 11520 14764 11572 14816
rect 13268 14764 13320 14816
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 2813 14662 2865 14714
rect 2877 14662 2929 14714
rect 2941 14662 2993 14714
rect 3005 14662 3057 14714
rect 3069 14662 3121 14714
rect 6539 14662 6591 14714
rect 6603 14662 6655 14714
rect 6667 14662 6719 14714
rect 6731 14662 6783 14714
rect 6795 14662 6847 14714
rect 10265 14662 10317 14714
rect 10329 14662 10381 14714
rect 10393 14662 10445 14714
rect 10457 14662 10509 14714
rect 10521 14662 10573 14714
rect 13991 14662 14043 14714
rect 14055 14662 14107 14714
rect 14119 14662 14171 14714
rect 14183 14662 14235 14714
rect 14247 14662 14299 14714
rect 4712 14560 4764 14612
rect 7288 14560 7340 14612
rect 7472 14560 7524 14612
rect 5540 14492 5592 14544
rect 6184 14492 6236 14544
rect 7380 14492 7432 14544
rect 5264 14399 5316 14408
rect 5264 14365 5273 14399
rect 5273 14365 5307 14399
rect 5307 14365 5316 14399
rect 5264 14356 5316 14365
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 7380 14356 7432 14408
rect 9128 14560 9180 14612
rect 9864 14560 9916 14612
rect 10048 14560 10100 14612
rect 12256 14603 12308 14612
rect 12256 14569 12265 14603
rect 12265 14569 12299 14603
rect 12299 14569 12308 14603
rect 12256 14560 12308 14569
rect 15292 14560 15344 14612
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 12992 14492 13044 14544
rect 8852 14424 8904 14476
rect 9496 14424 9548 14476
rect 9772 14424 9824 14476
rect 5724 14220 5776 14272
rect 5908 14220 5960 14272
rect 7012 14220 7064 14272
rect 7932 14263 7984 14272
rect 7932 14229 7941 14263
rect 7941 14229 7975 14263
rect 7975 14229 7984 14263
rect 7932 14220 7984 14229
rect 9404 14331 9456 14340
rect 9404 14297 9413 14331
rect 9413 14297 9447 14331
rect 9447 14297 9456 14331
rect 9404 14288 9456 14297
rect 10140 14288 10192 14340
rect 11520 14288 11572 14340
rect 12440 14399 12492 14408
rect 12440 14365 12449 14399
rect 12449 14365 12483 14399
rect 12483 14365 12492 14399
rect 12440 14356 12492 14365
rect 12992 14356 13044 14408
rect 13176 14356 13228 14408
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 13820 14424 13872 14476
rect 10048 14220 10100 14272
rect 10692 14220 10744 14272
rect 11336 14220 11388 14272
rect 12348 14220 12400 14272
rect 13636 14220 13688 14272
rect 13912 14220 13964 14272
rect 15016 14356 15068 14408
rect 3473 14118 3525 14170
rect 3537 14118 3589 14170
rect 3601 14118 3653 14170
rect 3665 14118 3717 14170
rect 3729 14118 3781 14170
rect 7199 14118 7251 14170
rect 7263 14118 7315 14170
rect 7327 14118 7379 14170
rect 7391 14118 7443 14170
rect 7455 14118 7507 14170
rect 10925 14118 10977 14170
rect 10989 14118 11041 14170
rect 11053 14118 11105 14170
rect 11117 14118 11169 14170
rect 11181 14118 11233 14170
rect 14651 14118 14703 14170
rect 14715 14118 14767 14170
rect 14779 14118 14831 14170
rect 14843 14118 14895 14170
rect 14907 14118 14959 14170
rect 4160 14016 4212 14068
rect 4804 14016 4856 14068
rect 5448 14059 5500 14068
rect 5448 14025 5457 14059
rect 5457 14025 5491 14059
rect 5491 14025 5500 14059
rect 5448 14016 5500 14025
rect 5724 14016 5776 14068
rect 7932 14016 7984 14068
rect 9404 14016 9456 14068
rect 9772 14016 9824 14068
rect 4988 13948 5040 14000
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 4620 13880 4672 13932
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 11428 14016 11480 14068
rect 11980 14016 12032 14068
rect 11520 13948 11572 14000
rect 10692 13880 10744 13932
rect 15568 14016 15620 14068
rect 14464 13948 14516 14000
rect 3884 13855 3936 13864
rect 3884 13821 3893 13855
rect 3893 13821 3927 13855
rect 3927 13821 3936 13855
rect 3884 13812 3936 13821
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 9128 13855 9180 13864
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 9128 13812 9180 13821
rect 11060 13812 11112 13864
rect 13084 13855 13136 13864
rect 13084 13821 13093 13855
rect 13093 13821 13127 13855
rect 13127 13821 13136 13855
rect 13084 13812 13136 13821
rect 15016 13812 15068 13864
rect 2504 13719 2556 13728
rect 2504 13685 2513 13719
rect 2513 13685 2547 13719
rect 2547 13685 2556 13719
rect 2504 13676 2556 13685
rect 14556 13676 14608 13728
rect 2813 13574 2865 13626
rect 2877 13574 2929 13626
rect 2941 13574 2993 13626
rect 3005 13574 3057 13626
rect 3069 13574 3121 13626
rect 6539 13574 6591 13626
rect 6603 13574 6655 13626
rect 6667 13574 6719 13626
rect 6731 13574 6783 13626
rect 6795 13574 6847 13626
rect 10265 13574 10317 13626
rect 10329 13574 10381 13626
rect 10393 13574 10445 13626
rect 10457 13574 10509 13626
rect 10521 13574 10573 13626
rect 13991 13574 14043 13626
rect 14055 13574 14107 13626
rect 14119 13574 14171 13626
rect 14183 13574 14235 13626
rect 14247 13574 14299 13626
rect 11060 13515 11112 13524
rect 11060 13481 11069 13515
rect 11069 13481 11103 13515
rect 11103 13481 11112 13515
rect 11060 13472 11112 13481
rect 13084 13472 13136 13524
rect 11336 13404 11388 13456
rect 2504 13336 2556 13388
rect 9680 13336 9732 13388
rect 10692 13336 10744 13388
rect 3148 13268 3200 13320
rect 3332 13268 3384 13320
rect 4344 13311 4396 13320
rect 4344 13277 4353 13311
rect 4353 13277 4387 13311
rect 4387 13277 4396 13311
rect 4344 13268 4396 13277
rect 6920 13268 6972 13320
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 7564 13200 7616 13252
rect 8300 13200 8352 13252
rect 10508 13311 10560 13320
rect 10508 13277 10517 13311
rect 10517 13277 10551 13311
rect 10551 13277 10560 13311
rect 10508 13268 10560 13277
rect 13636 13311 13688 13320
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 14556 13379 14608 13388
rect 14556 13345 14565 13379
rect 14565 13345 14599 13379
rect 14599 13345 14608 13379
rect 14556 13336 14608 13345
rect 13636 13268 13688 13277
rect 11428 13200 11480 13252
rect 13912 13200 13964 13252
rect 1952 13132 2004 13184
rect 3056 13132 3108 13184
rect 3884 13132 3936 13184
rect 9220 13175 9272 13184
rect 9220 13141 9229 13175
rect 9229 13141 9263 13175
rect 9263 13141 9272 13175
rect 9220 13132 9272 13141
rect 10600 13132 10652 13184
rect 13728 13132 13780 13184
rect 14556 13132 14608 13184
rect 3473 13030 3525 13082
rect 3537 13030 3589 13082
rect 3601 13030 3653 13082
rect 3665 13030 3717 13082
rect 3729 13030 3781 13082
rect 7199 13030 7251 13082
rect 7263 13030 7315 13082
rect 7327 13030 7379 13082
rect 7391 13030 7443 13082
rect 7455 13030 7507 13082
rect 10925 13030 10977 13082
rect 10989 13030 11041 13082
rect 11053 13030 11105 13082
rect 11117 13030 11169 13082
rect 11181 13030 11233 13082
rect 14651 13030 14703 13082
rect 14715 13030 14767 13082
rect 14779 13030 14831 13082
rect 14843 13030 14895 13082
rect 14907 13030 14959 13082
rect 3148 12928 3200 12980
rect 3424 12928 3476 12980
rect 2872 12860 2924 12912
rect 4988 12928 5040 12980
rect 7564 12928 7616 12980
rect 9036 12928 9088 12980
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 2136 12767 2188 12776
rect 2136 12733 2145 12767
rect 2145 12733 2179 12767
rect 2179 12733 2188 12767
rect 2136 12724 2188 12733
rect 2688 12724 2740 12776
rect 3884 12656 3936 12708
rect 4804 12835 4856 12844
rect 4804 12801 4813 12835
rect 4813 12801 4847 12835
rect 4847 12801 4856 12835
rect 4804 12792 4856 12801
rect 5080 12792 5132 12844
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5448 12835 5500 12844
rect 5448 12801 5457 12835
rect 5457 12801 5491 12835
rect 5491 12801 5500 12835
rect 5448 12792 5500 12801
rect 7104 12792 7156 12844
rect 9220 12928 9272 12980
rect 8392 12792 8444 12844
rect 10140 12860 10192 12912
rect 10600 12860 10652 12912
rect 10508 12792 10560 12844
rect 5908 12724 5960 12776
rect 6460 12724 6512 12776
rect 1952 12588 2004 12640
rect 2872 12588 2924 12640
rect 3148 12588 3200 12640
rect 6000 12656 6052 12708
rect 5540 12631 5592 12640
rect 5540 12597 5549 12631
rect 5549 12597 5583 12631
rect 5583 12597 5592 12631
rect 5540 12588 5592 12597
rect 8484 12631 8536 12640
rect 8484 12597 8493 12631
rect 8493 12597 8527 12631
rect 8527 12597 8536 12631
rect 8484 12588 8536 12597
rect 8852 12767 8904 12776
rect 8852 12733 8861 12767
rect 8861 12733 8895 12767
rect 8895 12733 8904 12767
rect 8852 12724 8904 12733
rect 9864 12588 9916 12640
rect 10140 12588 10192 12640
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 10692 12631 10744 12640
rect 10692 12597 10701 12631
rect 10701 12597 10735 12631
rect 10735 12597 10744 12631
rect 10692 12588 10744 12597
rect 12992 12792 13044 12844
rect 13452 12792 13504 12844
rect 14556 12792 14608 12844
rect 11152 12767 11204 12776
rect 11152 12733 11161 12767
rect 11161 12733 11195 12767
rect 11195 12733 11204 12767
rect 11152 12724 11204 12733
rect 11336 12656 11388 12708
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 10876 12588 10928 12640
rect 11612 12588 11664 12640
rect 12164 12631 12216 12640
rect 12164 12597 12173 12631
rect 12173 12597 12207 12631
rect 12207 12597 12216 12631
rect 12164 12588 12216 12597
rect 13360 12588 13412 12640
rect 13820 12631 13872 12640
rect 13820 12597 13829 12631
rect 13829 12597 13863 12631
rect 13863 12597 13872 12631
rect 13820 12588 13872 12597
rect 2813 12486 2865 12538
rect 2877 12486 2929 12538
rect 2941 12486 2993 12538
rect 3005 12486 3057 12538
rect 3069 12486 3121 12538
rect 6539 12486 6591 12538
rect 6603 12486 6655 12538
rect 6667 12486 6719 12538
rect 6731 12486 6783 12538
rect 6795 12486 6847 12538
rect 10265 12486 10317 12538
rect 10329 12486 10381 12538
rect 10393 12486 10445 12538
rect 10457 12486 10509 12538
rect 10521 12486 10573 12538
rect 13991 12486 14043 12538
rect 14055 12486 14107 12538
rect 14119 12486 14171 12538
rect 14183 12486 14235 12538
rect 14247 12486 14299 12538
rect 6552 12427 6604 12436
rect 6552 12393 6561 12427
rect 6561 12393 6595 12427
rect 6595 12393 6604 12427
rect 6552 12384 6604 12393
rect 9864 12384 9916 12436
rect 7012 12316 7064 12368
rect 3884 12248 3936 12300
rect 5172 12180 5224 12232
rect 5264 12223 5316 12232
rect 5264 12189 5273 12223
rect 5273 12189 5307 12223
rect 5307 12189 5316 12223
rect 5264 12180 5316 12189
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 8116 12248 8168 12300
rect 9772 12248 9824 12300
rect 10140 12248 10192 12300
rect 1952 12044 2004 12096
rect 3424 12112 3476 12164
rect 3976 12112 4028 12164
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 7656 12180 7708 12189
rect 7748 12155 7800 12164
rect 7748 12121 7757 12155
rect 7757 12121 7791 12155
rect 7791 12121 7800 12155
rect 7748 12112 7800 12121
rect 8484 12223 8536 12232
rect 8484 12189 8493 12223
rect 8493 12189 8527 12223
rect 8527 12189 8536 12223
rect 8484 12180 8536 12189
rect 9128 12180 9180 12232
rect 9680 12180 9732 12232
rect 10784 12291 10836 12300
rect 10784 12257 10793 12291
rect 10793 12257 10827 12291
rect 10827 12257 10836 12291
rect 10784 12248 10836 12257
rect 4528 12044 4580 12096
rect 4620 12087 4672 12096
rect 4620 12053 4629 12087
rect 4629 12053 4663 12087
rect 4663 12053 4672 12087
rect 4620 12044 4672 12053
rect 4712 12087 4764 12096
rect 4712 12053 4721 12087
rect 4721 12053 4755 12087
rect 4755 12053 4764 12087
rect 4712 12044 4764 12053
rect 5080 12044 5132 12096
rect 6736 12044 6788 12096
rect 10600 12112 10652 12164
rect 8208 12044 8260 12096
rect 8576 12044 8628 12096
rect 10876 12180 10928 12232
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 11704 12384 11756 12436
rect 12164 12384 12216 12436
rect 12808 12316 12860 12368
rect 11980 12248 12032 12300
rect 12716 12180 12768 12232
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 13544 12180 13596 12232
rect 14556 12180 14608 12232
rect 10784 12044 10836 12096
rect 11704 12112 11756 12164
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 13820 12044 13872 12096
rect 3473 11942 3525 11994
rect 3537 11942 3589 11994
rect 3601 11942 3653 11994
rect 3665 11942 3717 11994
rect 3729 11942 3781 11994
rect 7199 11942 7251 11994
rect 7263 11942 7315 11994
rect 7327 11942 7379 11994
rect 7391 11942 7443 11994
rect 7455 11942 7507 11994
rect 10925 11942 10977 11994
rect 10989 11942 11041 11994
rect 11053 11942 11105 11994
rect 11117 11942 11169 11994
rect 11181 11942 11233 11994
rect 14651 11942 14703 11994
rect 14715 11942 14767 11994
rect 14779 11942 14831 11994
rect 14843 11942 14895 11994
rect 14907 11942 14959 11994
rect 2136 11840 2188 11892
rect 3884 11840 3936 11892
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 7748 11840 7800 11892
rect 3240 11772 3292 11824
rect 3516 11772 3568 11824
rect 2688 11704 2740 11756
rect 3332 11704 3384 11756
rect 3976 11772 4028 11824
rect 4436 11747 4488 11756
rect 3240 11679 3292 11688
rect 3240 11645 3249 11679
rect 3249 11645 3283 11679
rect 3283 11645 3292 11679
rect 3240 11636 3292 11645
rect 4436 11713 4445 11747
rect 4445 11713 4479 11747
rect 4479 11713 4488 11747
rect 4436 11704 4488 11713
rect 1952 11568 2004 11620
rect 4252 11636 4304 11688
rect 4344 11636 4396 11688
rect 4712 11679 4764 11688
rect 4712 11645 4721 11679
rect 4721 11645 4755 11679
rect 4755 11645 4764 11679
rect 4712 11636 4764 11645
rect 5448 11636 5500 11688
rect 6828 11772 6880 11824
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 8484 11840 8536 11892
rect 10140 11840 10192 11892
rect 13176 11840 13228 11892
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 3516 11611 3568 11620
rect 3516 11577 3525 11611
rect 3525 11577 3559 11611
rect 3559 11577 3568 11611
rect 3516 11568 3568 11577
rect 3792 11568 3844 11620
rect 8024 11636 8076 11688
rect 11704 11636 11756 11688
rect 3148 11500 3200 11552
rect 3884 11500 3936 11552
rect 4068 11500 4120 11552
rect 8576 11611 8628 11620
rect 8576 11577 8585 11611
rect 8585 11577 8619 11611
rect 8619 11577 8628 11611
rect 8576 11568 8628 11577
rect 11612 11611 11664 11620
rect 11612 11577 11621 11611
rect 11621 11577 11655 11611
rect 11655 11577 11664 11611
rect 11612 11568 11664 11577
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 8484 11500 8536 11552
rect 11980 11704 12032 11756
rect 12808 11747 12860 11756
rect 12808 11713 12817 11747
rect 12817 11713 12851 11747
rect 12851 11713 12860 11747
rect 12808 11704 12860 11713
rect 14372 11704 14424 11756
rect 14556 11679 14608 11688
rect 14556 11645 14565 11679
rect 14565 11645 14599 11679
rect 14599 11645 14608 11679
rect 14556 11636 14608 11645
rect 13544 11500 13596 11552
rect 2813 11398 2865 11450
rect 2877 11398 2929 11450
rect 2941 11398 2993 11450
rect 3005 11398 3057 11450
rect 3069 11398 3121 11450
rect 6539 11398 6591 11450
rect 6603 11398 6655 11450
rect 6667 11398 6719 11450
rect 6731 11398 6783 11450
rect 6795 11398 6847 11450
rect 10265 11398 10317 11450
rect 10329 11398 10381 11450
rect 10393 11398 10445 11450
rect 10457 11398 10509 11450
rect 10521 11398 10573 11450
rect 13991 11398 14043 11450
rect 14055 11398 14107 11450
rect 14119 11398 14171 11450
rect 14183 11398 14235 11450
rect 14247 11398 14299 11450
rect 3332 11296 3384 11348
rect 3240 11228 3292 11280
rect 4160 11296 4212 11348
rect 4252 11339 4304 11348
rect 4252 11305 4261 11339
rect 4261 11305 4295 11339
rect 4295 11305 4304 11339
rect 4252 11296 4304 11305
rect 4344 11296 4396 11348
rect 4436 11296 4488 11348
rect 4528 11339 4580 11348
rect 4528 11305 4537 11339
rect 4537 11305 4571 11339
rect 4571 11305 4580 11339
rect 4528 11296 4580 11305
rect 5264 11296 5316 11348
rect 5540 11296 5592 11348
rect 7564 11296 7616 11348
rect 8116 11296 8168 11348
rect 8208 11296 8260 11348
rect 3976 11228 4028 11280
rect 3240 11024 3292 11076
rect 2780 10956 2832 11008
rect 2964 10956 3016 11008
rect 4068 11203 4120 11220
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11168 4120 11169
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 7012 11228 7064 11280
rect 8024 11271 8076 11280
rect 8024 11237 8033 11271
rect 8033 11237 8067 11271
rect 8067 11237 8076 11271
rect 8024 11228 8076 11237
rect 5540 11160 5592 11212
rect 6000 11160 6052 11212
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 5080 11135 5132 11144
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 7748 11160 7800 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 11336 11160 11388 11212
rect 11796 11203 11848 11212
rect 11796 11169 11805 11203
rect 11805 11169 11839 11203
rect 11839 11169 11848 11203
rect 11796 11160 11848 11169
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 11520 11092 11572 11144
rect 12716 11228 12768 11280
rect 13452 11228 13504 11280
rect 13544 11228 13596 11280
rect 12624 11160 12676 11212
rect 8484 11024 8536 11076
rect 4252 10956 4304 11008
rect 5356 10956 5408 11008
rect 7656 10956 7708 11008
rect 10600 10956 10652 11008
rect 11428 10956 11480 11008
rect 13360 11092 13412 11144
rect 13728 11160 13780 11212
rect 15016 11092 15068 11144
rect 13728 11024 13780 11076
rect 12348 10956 12400 11008
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12440 10956 12492 10965
rect 12532 10999 12584 11008
rect 12532 10965 12541 10999
rect 12541 10965 12575 10999
rect 12575 10965 12584 10999
rect 12532 10956 12584 10965
rect 14372 11024 14424 11076
rect 15384 11024 15436 11076
rect 14464 10956 14516 11008
rect 14556 10956 14608 11008
rect 3473 10854 3525 10906
rect 3537 10854 3589 10906
rect 3601 10854 3653 10906
rect 3665 10854 3717 10906
rect 3729 10854 3781 10906
rect 7199 10854 7251 10906
rect 7263 10854 7315 10906
rect 7327 10854 7379 10906
rect 7391 10854 7443 10906
rect 7455 10854 7507 10906
rect 10925 10854 10977 10906
rect 10989 10854 11041 10906
rect 11053 10854 11105 10906
rect 11117 10854 11169 10906
rect 11181 10854 11233 10906
rect 14651 10854 14703 10906
rect 14715 10854 14767 10906
rect 14779 10854 14831 10906
rect 14843 10854 14895 10906
rect 14907 10854 14959 10906
rect 3148 10752 3200 10804
rect 9496 10752 9548 10804
rect 9680 10752 9732 10804
rect 10784 10752 10836 10804
rect 11336 10752 11388 10804
rect 11612 10752 11664 10804
rect 12808 10752 12860 10804
rect 2872 10684 2924 10736
rect 8484 10684 8536 10736
rect 14372 10684 14424 10736
rect 14556 10684 14608 10736
rect 940 10616 992 10668
rect 4160 10616 4212 10668
rect 4988 10659 5040 10668
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 5356 10616 5408 10668
rect 5540 10616 5592 10668
rect 9220 10616 9272 10668
rect 9588 10659 9640 10668
rect 9588 10625 9597 10659
rect 9597 10625 9631 10659
rect 9631 10625 9640 10659
rect 9588 10616 9640 10625
rect 11428 10616 11480 10668
rect 11796 10616 11848 10668
rect 13636 10616 13688 10668
rect 15016 10795 15068 10804
rect 15016 10761 15025 10795
rect 15025 10761 15059 10795
rect 15059 10761 15068 10795
rect 15016 10752 15068 10761
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 2228 10591 2280 10600
rect 2228 10557 2237 10591
rect 2237 10557 2271 10591
rect 2271 10557 2280 10591
rect 2228 10548 2280 10557
rect 2964 10548 3016 10600
rect 4620 10591 4672 10600
rect 4620 10557 4629 10591
rect 4629 10557 4663 10591
rect 4663 10557 4672 10591
rect 4620 10548 4672 10557
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 12440 10548 12492 10600
rect 15108 10548 15160 10600
rect 12624 10480 12676 10532
rect 3792 10455 3844 10464
rect 3792 10421 3801 10455
rect 3801 10421 3835 10455
rect 3835 10421 3844 10455
rect 3792 10412 3844 10421
rect 5172 10412 5224 10464
rect 11704 10412 11756 10464
rect 12348 10455 12400 10464
rect 12348 10421 12357 10455
rect 12357 10421 12391 10455
rect 12391 10421 12400 10455
rect 12348 10412 12400 10421
rect 2813 10310 2865 10362
rect 2877 10310 2929 10362
rect 2941 10310 2993 10362
rect 3005 10310 3057 10362
rect 3069 10310 3121 10362
rect 6539 10310 6591 10362
rect 6603 10310 6655 10362
rect 6667 10310 6719 10362
rect 6731 10310 6783 10362
rect 6795 10310 6847 10362
rect 10265 10310 10317 10362
rect 10329 10310 10381 10362
rect 10393 10310 10445 10362
rect 10457 10310 10509 10362
rect 10521 10310 10573 10362
rect 13991 10310 14043 10362
rect 14055 10310 14107 10362
rect 14119 10310 14171 10362
rect 14183 10310 14235 10362
rect 14247 10310 14299 10362
rect 2228 10208 2280 10260
rect 3792 10208 3844 10260
rect 5540 10251 5592 10260
rect 5540 10217 5549 10251
rect 5549 10217 5583 10251
rect 5583 10217 5592 10251
rect 5540 10208 5592 10217
rect 7104 10251 7156 10260
rect 7104 10217 7113 10251
rect 7113 10217 7147 10251
rect 7147 10217 7156 10251
rect 7104 10208 7156 10217
rect 7196 10208 7248 10260
rect 12624 10208 12676 10260
rect 15016 10208 15068 10260
rect 3148 10072 3200 10124
rect 2780 10004 2832 10056
rect 13728 10140 13780 10192
rect 7656 10115 7708 10124
rect 7656 10081 7665 10115
rect 7665 10081 7699 10115
rect 7699 10081 7708 10115
rect 7656 10072 7708 10081
rect 3884 10004 3936 10056
rect 9680 10072 9732 10124
rect 11336 10072 11388 10124
rect 13636 10072 13688 10124
rect 13912 10072 13964 10124
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 4068 9936 4120 9988
rect 6920 9936 6972 9988
rect 9588 9936 9640 9988
rect 11520 9936 11572 9988
rect 3240 9868 3292 9920
rect 4160 9868 4212 9920
rect 15016 9868 15068 9920
rect 3473 9766 3525 9818
rect 3537 9766 3589 9818
rect 3601 9766 3653 9818
rect 3665 9766 3717 9818
rect 3729 9766 3781 9818
rect 7199 9766 7251 9818
rect 7263 9766 7315 9818
rect 7327 9766 7379 9818
rect 7391 9766 7443 9818
rect 7455 9766 7507 9818
rect 10925 9766 10977 9818
rect 10989 9766 11041 9818
rect 11053 9766 11105 9818
rect 11117 9766 11169 9818
rect 11181 9766 11233 9818
rect 14651 9766 14703 9818
rect 14715 9766 14767 9818
rect 14779 9766 14831 9818
rect 14843 9766 14895 9818
rect 14907 9766 14959 9818
rect 4160 9664 4212 9716
rect 11336 9664 11388 9716
rect 12256 9664 12308 9716
rect 12624 9664 12676 9716
rect 15108 9707 15160 9716
rect 15108 9673 15117 9707
rect 15117 9673 15151 9707
rect 15151 9673 15160 9707
rect 15108 9664 15160 9673
rect 3148 9596 3200 9648
rect 13912 9596 13964 9648
rect 14372 9596 14424 9648
rect 3332 9528 3384 9580
rect 3884 9571 3936 9580
rect 3884 9537 3893 9571
rect 3893 9537 3927 9571
rect 3927 9537 3936 9571
rect 3884 9528 3936 9537
rect 3976 9528 4028 9580
rect 4068 9528 4120 9580
rect 4620 9460 4672 9512
rect 4804 9503 4856 9512
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 5172 9571 5224 9580
rect 5172 9537 5181 9571
rect 5181 9537 5215 9571
rect 5215 9537 5224 9571
rect 5172 9528 5224 9537
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 10784 9528 10836 9580
rect 11336 9528 11388 9580
rect 9220 9460 9272 9512
rect 11704 9460 11756 9512
rect 12256 9460 12308 9512
rect 12808 9528 12860 9580
rect 12532 9460 12584 9512
rect 2688 9324 2740 9376
rect 3792 9324 3844 9376
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 4896 9367 4948 9376
rect 4896 9333 4905 9367
rect 4905 9333 4939 9367
rect 4939 9333 4948 9367
rect 4896 9324 4948 9333
rect 9680 9324 9732 9376
rect 10600 9324 10652 9376
rect 11520 9324 11572 9376
rect 11704 9324 11756 9376
rect 11888 9324 11940 9376
rect 15384 9324 15436 9376
rect 2813 9222 2865 9274
rect 2877 9222 2929 9274
rect 2941 9222 2993 9274
rect 3005 9222 3057 9274
rect 3069 9222 3121 9274
rect 6539 9222 6591 9274
rect 6603 9222 6655 9274
rect 6667 9222 6719 9274
rect 6731 9222 6783 9274
rect 6795 9222 6847 9274
rect 10265 9222 10317 9274
rect 10329 9222 10381 9274
rect 10393 9222 10445 9274
rect 10457 9222 10509 9274
rect 10521 9222 10573 9274
rect 13991 9222 14043 9274
rect 14055 9222 14107 9274
rect 14119 9222 14171 9274
rect 14183 9222 14235 9274
rect 14247 9222 14299 9274
rect 4068 9120 4120 9172
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 4804 9120 4856 9172
rect 8208 9120 8260 9172
rect 11152 9120 11204 9172
rect 5448 9052 5500 9104
rect 7196 9052 7248 9104
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 3240 8916 3292 8968
rect 3056 8780 3108 8832
rect 4528 8916 4580 8968
rect 8208 8984 8260 9036
rect 7196 8916 7248 8968
rect 8024 8959 8076 8968
rect 8024 8925 8033 8959
rect 8033 8925 8067 8959
rect 8067 8925 8076 8959
rect 8024 8916 8076 8925
rect 8116 8916 8168 8968
rect 8576 9052 8628 9104
rect 11520 9052 11572 9104
rect 11612 9052 11664 9104
rect 12256 9095 12308 9104
rect 12256 9061 12265 9095
rect 12265 9061 12299 9095
rect 12299 9061 12308 9095
rect 12256 9052 12308 9061
rect 12440 9052 12492 9104
rect 15016 9120 15068 9172
rect 15384 9120 15436 9172
rect 11244 9027 11296 9036
rect 11244 8993 11253 9027
rect 11253 8993 11287 9027
rect 11287 8993 11296 9027
rect 11244 8984 11296 8993
rect 14464 8984 14516 9036
rect 7012 8848 7064 8900
rect 9588 8916 9640 8968
rect 9772 8848 9824 8900
rect 7932 8780 7984 8832
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 8760 8780 8812 8832
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 10232 8823 10284 8832
rect 10232 8789 10241 8823
rect 10241 8789 10275 8823
rect 10275 8789 10284 8823
rect 10232 8780 10284 8789
rect 11152 8953 11204 8968
rect 11152 8919 11161 8953
rect 11161 8919 11195 8953
rect 11195 8919 11204 8953
rect 11152 8916 11204 8919
rect 11336 8848 11388 8900
rect 11704 8916 11756 8968
rect 11980 8916 12032 8968
rect 11888 8848 11940 8900
rect 14924 8984 14976 9036
rect 12440 8891 12492 8900
rect 12440 8857 12449 8891
rect 12449 8857 12483 8891
rect 12483 8857 12492 8891
rect 12440 8848 12492 8857
rect 13820 8848 13872 8900
rect 16028 8848 16080 8900
rect 12164 8780 12216 8832
rect 12624 8823 12676 8832
rect 12624 8789 12633 8823
rect 12633 8789 12667 8823
rect 12667 8789 12676 8823
rect 12624 8780 12676 8789
rect 14280 8780 14332 8832
rect 14740 8780 14792 8832
rect 15016 8780 15068 8832
rect 3473 8678 3525 8730
rect 3537 8678 3589 8730
rect 3601 8678 3653 8730
rect 3665 8678 3717 8730
rect 3729 8678 3781 8730
rect 7199 8678 7251 8730
rect 7263 8678 7315 8730
rect 7327 8678 7379 8730
rect 7391 8678 7443 8730
rect 7455 8678 7507 8730
rect 10925 8678 10977 8730
rect 10989 8678 11041 8730
rect 11053 8678 11105 8730
rect 11117 8678 11169 8730
rect 11181 8678 11233 8730
rect 14651 8678 14703 8730
rect 14715 8678 14767 8730
rect 14779 8678 14831 8730
rect 14843 8678 14895 8730
rect 14907 8678 14959 8730
rect 1860 8440 1912 8492
rect 4436 8576 4488 8628
rect 4528 8619 4580 8628
rect 4528 8585 4537 8619
rect 4537 8585 4571 8619
rect 4571 8585 4580 8619
rect 4528 8576 4580 8585
rect 3056 8508 3108 8560
rect 7288 8576 7340 8628
rect 9588 8576 9640 8628
rect 9220 8508 9272 8560
rect 4896 8440 4948 8492
rect 6276 8440 6328 8492
rect 9772 8508 9824 8560
rect 10232 8576 10284 8628
rect 12164 8619 12216 8628
rect 12164 8585 12173 8619
rect 12173 8585 12207 8619
rect 12207 8585 12216 8619
rect 12164 8576 12216 8585
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 13452 8508 13504 8560
rect 15384 8508 15436 8560
rect 6092 8372 6144 8424
rect 7104 8372 7156 8424
rect 3240 8236 3292 8288
rect 4804 8304 4856 8356
rect 10876 8440 10928 8492
rect 12624 8440 12676 8492
rect 8944 8372 8996 8424
rect 11060 8372 11112 8424
rect 11520 8415 11572 8424
rect 11520 8381 11529 8415
rect 11529 8381 11563 8415
rect 11563 8381 11572 8415
rect 11520 8372 11572 8381
rect 12716 8415 12768 8424
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 13452 8372 13504 8424
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 8116 8279 8168 8288
rect 8116 8245 8125 8279
rect 8125 8245 8159 8279
rect 8159 8245 8168 8279
rect 8116 8236 8168 8245
rect 10968 8236 11020 8288
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 2813 8134 2865 8186
rect 2877 8134 2929 8186
rect 2941 8134 2993 8186
rect 3005 8134 3057 8186
rect 3069 8134 3121 8186
rect 6539 8134 6591 8186
rect 6603 8134 6655 8186
rect 6667 8134 6719 8186
rect 6731 8134 6783 8186
rect 6795 8134 6847 8186
rect 10265 8134 10317 8186
rect 10329 8134 10381 8186
rect 10393 8134 10445 8186
rect 10457 8134 10509 8186
rect 10521 8134 10573 8186
rect 13991 8134 14043 8186
rect 14055 8134 14107 8186
rect 14119 8134 14171 8186
rect 14183 8134 14235 8186
rect 14247 8134 14299 8186
rect 3976 8032 4028 8084
rect 4436 8032 4488 8084
rect 8024 8032 8076 8084
rect 8760 8032 8812 8084
rect 11520 8032 11572 8084
rect 12256 8032 12308 8084
rect 11060 8007 11112 8016
rect 11060 7973 11069 8007
rect 11069 7973 11103 8007
rect 11103 7973 11112 8007
rect 11060 7964 11112 7973
rect 6276 7939 6328 7948
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3332 7828 3384 7837
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 7012 7896 7064 7948
rect 7288 7896 7340 7948
rect 7748 7896 7800 7948
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 5448 7828 5500 7880
rect 7932 7828 7984 7880
rect 8392 7871 8444 7880
rect 8392 7837 8401 7871
rect 8401 7837 8435 7871
rect 8435 7837 8444 7871
rect 8392 7828 8444 7837
rect 8944 7939 8996 7948
rect 8944 7905 8953 7939
rect 8953 7905 8987 7939
rect 8987 7905 8996 7939
rect 8944 7896 8996 7905
rect 9680 7896 9732 7948
rect 11336 7939 11388 7948
rect 11336 7905 11345 7939
rect 11345 7905 11379 7939
rect 11379 7905 11388 7939
rect 14372 7964 14424 8016
rect 11336 7896 11388 7905
rect 13820 7896 13872 7948
rect 14464 7896 14516 7948
rect 15108 7896 15160 7948
rect 3332 7692 3384 7744
rect 3976 7692 4028 7744
rect 4344 7735 4396 7744
rect 4344 7701 4353 7735
rect 4353 7701 4387 7735
rect 4387 7701 4396 7735
rect 4344 7692 4396 7701
rect 6828 7760 6880 7812
rect 7288 7760 7340 7812
rect 6920 7692 6972 7744
rect 8300 7760 8352 7812
rect 10968 7828 11020 7880
rect 11612 7828 11664 7880
rect 9220 7760 9272 7812
rect 13452 7828 13504 7880
rect 15200 7828 15252 7880
rect 12716 7760 12768 7812
rect 10784 7692 10836 7744
rect 14372 7692 14424 7744
rect 15292 7692 15344 7744
rect 3473 7590 3525 7642
rect 3537 7590 3589 7642
rect 3601 7590 3653 7642
rect 3665 7590 3717 7642
rect 3729 7590 3781 7642
rect 7199 7590 7251 7642
rect 7263 7590 7315 7642
rect 7327 7590 7379 7642
rect 7391 7590 7443 7642
rect 7455 7590 7507 7642
rect 10925 7590 10977 7642
rect 10989 7590 11041 7642
rect 11053 7590 11105 7642
rect 11117 7590 11169 7642
rect 11181 7590 11233 7642
rect 14651 7590 14703 7642
rect 14715 7590 14767 7642
rect 14779 7590 14831 7642
rect 14843 7590 14895 7642
rect 14907 7590 14959 7642
rect 3240 7488 3292 7540
rect 1860 7352 1912 7404
rect 4252 7488 4304 7540
rect 4344 7488 4396 7540
rect 5448 7488 5500 7540
rect 6000 7488 6052 7540
rect 3884 7352 3936 7404
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 7012 7420 7064 7472
rect 7748 7420 7800 7472
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 4160 7327 4212 7336
rect 4160 7293 4169 7327
rect 4169 7293 4203 7327
rect 4203 7293 4212 7327
rect 4160 7284 4212 7293
rect 4988 7284 5040 7336
rect 5264 7284 5316 7336
rect 4896 7216 4948 7268
rect 6276 7352 6328 7404
rect 7196 7284 7248 7336
rect 8208 7531 8260 7540
rect 8208 7497 8217 7531
rect 8217 7497 8251 7531
rect 8251 7497 8260 7531
rect 8208 7488 8260 7497
rect 8392 7488 8444 7540
rect 11336 7488 11388 7540
rect 12716 7488 12768 7540
rect 8576 7420 8628 7472
rect 9220 7352 9272 7404
rect 13452 7420 13504 7472
rect 14372 7420 14424 7472
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 15108 7488 15160 7540
rect 15200 7420 15252 7472
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 12440 7284 12492 7336
rect 14924 7284 14976 7336
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 3424 7148 3476 7200
rect 4252 7148 4304 7200
rect 6000 7148 6052 7200
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 9680 7216 9732 7268
rect 15108 7216 15160 7268
rect 8116 7148 8168 7200
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 9312 7191 9364 7200
rect 9312 7157 9321 7191
rect 9321 7157 9355 7191
rect 9355 7157 9364 7191
rect 9312 7148 9364 7157
rect 2813 7046 2865 7098
rect 2877 7046 2929 7098
rect 2941 7046 2993 7098
rect 3005 7046 3057 7098
rect 3069 7046 3121 7098
rect 6539 7046 6591 7098
rect 6603 7046 6655 7098
rect 6667 7046 6719 7098
rect 6731 7046 6783 7098
rect 6795 7046 6847 7098
rect 10265 7046 10317 7098
rect 10329 7046 10381 7098
rect 10393 7046 10445 7098
rect 10457 7046 10509 7098
rect 10521 7046 10573 7098
rect 13991 7046 14043 7098
rect 14055 7046 14107 7098
rect 14119 7046 14171 7098
rect 14183 7046 14235 7098
rect 14247 7046 14299 7098
rect 4160 6944 4212 6996
rect 4896 6987 4948 6996
rect 4896 6953 4905 6987
rect 4905 6953 4939 6987
rect 4939 6953 4948 6987
rect 4896 6944 4948 6953
rect 5080 6944 5132 6996
rect 7196 6944 7248 6996
rect 8208 6944 8260 6996
rect 11520 6944 11572 6996
rect 11704 6944 11756 6996
rect 13820 6944 13872 6996
rect 4068 6876 4120 6928
rect 5264 6876 5316 6928
rect 6736 6876 6788 6928
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 3240 6740 3292 6792
rect 3056 6604 3108 6656
rect 3976 6604 4028 6656
rect 4252 6740 4304 6792
rect 5448 6808 5500 6860
rect 7104 6808 7156 6860
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 6184 6740 6236 6792
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7288 6783 7340 6792
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 7932 6808 7984 6860
rect 8576 6808 8628 6860
rect 12716 6876 12768 6928
rect 4436 6672 4488 6724
rect 6092 6672 6144 6724
rect 7012 6672 7064 6724
rect 8392 6740 8444 6792
rect 12072 6740 12124 6792
rect 13912 6740 13964 6792
rect 14372 6808 14424 6860
rect 14464 6740 14516 6792
rect 14924 6740 14976 6792
rect 8300 6672 8352 6724
rect 10784 6672 10836 6724
rect 13452 6672 13504 6724
rect 12164 6647 12216 6656
rect 12164 6613 12173 6647
rect 12173 6613 12207 6647
rect 12207 6613 12216 6647
rect 12164 6604 12216 6613
rect 15108 6672 15160 6724
rect 14556 6604 14608 6656
rect 3473 6502 3525 6554
rect 3537 6502 3589 6554
rect 3601 6502 3653 6554
rect 3665 6502 3717 6554
rect 3729 6502 3781 6554
rect 7199 6502 7251 6554
rect 7263 6502 7315 6554
rect 7327 6502 7379 6554
rect 7391 6502 7443 6554
rect 7455 6502 7507 6554
rect 10925 6502 10977 6554
rect 10989 6502 11041 6554
rect 11053 6502 11105 6554
rect 11117 6502 11169 6554
rect 11181 6502 11233 6554
rect 14651 6502 14703 6554
rect 14715 6502 14767 6554
rect 14779 6502 14831 6554
rect 14843 6502 14895 6554
rect 14907 6502 14959 6554
rect 3884 6400 3936 6452
rect 4160 6400 4212 6452
rect 7104 6400 7156 6452
rect 8300 6400 8352 6452
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 12164 6400 12216 6452
rect 3240 6332 3292 6384
rect 3148 6264 3200 6316
rect 3332 6264 3384 6316
rect 4068 6264 4120 6316
rect 4436 6264 4488 6316
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 5080 6264 5132 6316
rect 5172 6264 5224 6316
rect 5448 6264 5500 6316
rect 8944 6264 8996 6316
rect 10876 6264 10928 6316
rect 11888 6264 11940 6316
rect 12072 6264 12124 6316
rect 3976 6196 4028 6205
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 5632 6128 5684 6180
rect 11704 6128 11756 6180
rect 12348 6128 12400 6180
rect 7104 6060 7156 6112
rect 2813 5958 2865 6010
rect 2877 5958 2929 6010
rect 2941 5958 2993 6010
rect 3005 5958 3057 6010
rect 3069 5958 3121 6010
rect 6539 5958 6591 6010
rect 6603 5958 6655 6010
rect 6667 5958 6719 6010
rect 6731 5958 6783 6010
rect 6795 5958 6847 6010
rect 10265 5958 10317 6010
rect 10329 5958 10381 6010
rect 10393 5958 10445 6010
rect 10457 5958 10509 6010
rect 10521 5958 10573 6010
rect 13991 5958 14043 6010
rect 14055 5958 14107 6010
rect 14119 5958 14171 6010
rect 14183 5958 14235 6010
rect 14247 5958 14299 6010
rect 4436 5856 4488 5908
rect 9864 5856 9916 5908
rect 4712 5788 4764 5840
rect 12624 5788 12676 5840
rect 14372 5788 14424 5840
rect 2688 5652 2740 5704
rect 2780 5584 2832 5636
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 5540 5720 5592 5772
rect 3976 5652 4028 5704
rect 3148 5516 3200 5568
rect 3884 5627 3936 5636
rect 3884 5593 3893 5627
rect 3893 5593 3927 5627
rect 3927 5593 3936 5627
rect 3884 5584 3936 5593
rect 4068 5627 4120 5636
rect 4068 5593 4077 5627
rect 4077 5593 4111 5627
rect 4111 5593 4120 5627
rect 4068 5584 4120 5593
rect 6460 5652 6512 5704
rect 7012 5652 7064 5704
rect 10600 5652 10652 5704
rect 11980 5652 12032 5704
rect 12900 5720 12952 5772
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 13912 5652 13964 5704
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 11520 5584 11572 5636
rect 12440 5584 12492 5636
rect 6184 5516 6236 5568
rect 6828 5559 6880 5568
rect 6828 5525 6837 5559
rect 6837 5525 6871 5559
rect 6871 5525 6880 5559
rect 6828 5516 6880 5525
rect 8300 5516 8352 5568
rect 8576 5516 8628 5568
rect 8944 5516 8996 5568
rect 12716 5516 12768 5568
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 3473 5414 3525 5466
rect 3537 5414 3589 5466
rect 3601 5414 3653 5466
rect 3665 5414 3717 5466
rect 3729 5414 3781 5466
rect 7199 5414 7251 5466
rect 7263 5414 7315 5466
rect 7327 5414 7379 5466
rect 7391 5414 7443 5466
rect 7455 5414 7507 5466
rect 10925 5414 10977 5466
rect 10989 5414 11041 5466
rect 11053 5414 11105 5466
rect 11117 5414 11169 5466
rect 11181 5414 11233 5466
rect 14651 5414 14703 5466
rect 14715 5414 14767 5466
rect 14779 5414 14831 5466
rect 14843 5414 14895 5466
rect 14907 5414 14959 5466
rect 3332 5312 3384 5364
rect 3976 5244 4028 5296
rect 4620 5312 4672 5364
rect 7564 5312 7616 5364
rect 6092 5287 6144 5296
rect 6092 5253 6101 5287
rect 6101 5253 6135 5287
rect 6135 5253 6144 5287
rect 6092 5244 6144 5253
rect 3056 5176 3108 5228
rect 3424 5176 3476 5228
rect 3884 5176 3936 5228
rect 4988 5176 5040 5228
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 3332 5108 3384 5160
rect 3792 5151 3844 5160
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 4068 5108 4120 5160
rect 4896 5108 4948 5160
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 9312 5176 9364 5228
rect 5172 5040 5224 5092
rect 5448 5040 5500 5092
rect 2504 4972 2556 5024
rect 3240 4972 3292 5024
rect 4068 4972 4120 5024
rect 4620 5015 4672 5024
rect 4620 4981 4629 5015
rect 4629 4981 4663 5015
rect 4663 4981 4672 5015
rect 4620 4972 4672 4981
rect 6000 4972 6052 5024
rect 6828 4972 6880 5024
rect 7656 5040 7708 5092
rect 7564 4972 7616 5024
rect 9128 4972 9180 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 11520 5355 11572 5364
rect 11520 5321 11529 5355
rect 11529 5321 11563 5355
rect 11563 5321 11572 5355
rect 11520 5312 11572 5321
rect 12348 5244 12400 5296
rect 10600 5176 10652 5228
rect 11520 5176 11572 5228
rect 12716 5312 12768 5364
rect 13452 5312 13504 5364
rect 13728 5312 13780 5364
rect 9864 5151 9916 5160
rect 9864 5117 9873 5151
rect 9873 5117 9907 5151
rect 9907 5117 9916 5151
rect 9864 5108 9916 5117
rect 10692 5151 10744 5160
rect 10692 5117 10701 5151
rect 10701 5117 10735 5151
rect 10735 5117 10744 5151
rect 10692 5108 10744 5117
rect 9956 5040 10008 5092
rect 11428 5040 11480 5092
rect 12072 5151 12124 5160
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 12624 5176 12676 5228
rect 12808 5219 12860 5228
rect 12808 5185 12817 5219
rect 12817 5185 12851 5219
rect 12851 5185 12860 5219
rect 12808 5176 12860 5185
rect 12900 5176 12952 5228
rect 14096 5244 14148 5296
rect 15384 5312 15436 5364
rect 10968 4972 11020 5024
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 12072 4972 12124 5024
rect 12532 4972 12584 5024
rect 2813 4870 2865 4922
rect 2877 4870 2929 4922
rect 2941 4870 2993 4922
rect 3005 4870 3057 4922
rect 3069 4870 3121 4922
rect 6539 4870 6591 4922
rect 6603 4870 6655 4922
rect 6667 4870 6719 4922
rect 6731 4870 6783 4922
rect 6795 4870 6847 4922
rect 10265 4870 10317 4922
rect 10329 4870 10381 4922
rect 10393 4870 10445 4922
rect 10457 4870 10509 4922
rect 10521 4870 10573 4922
rect 13991 4870 14043 4922
rect 14055 4870 14107 4922
rect 14119 4870 14171 4922
rect 14183 4870 14235 4922
rect 14247 4870 14299 4922
rect 3792 4768 3844 4820
rect 4344 4768 4396 4820
rect 4620 4768 4672 4820
rect 4896 4768 4948 4820
rect 5172 4768 5224 4820
rect 6000 4768 6052 4820
rect 6092 4768 6144 4820
rect 7196 4768 7248 4820
rect 1860 4675 1912 4684
rect 1860 4641 1869 4675
rect 1869 4641 1903 4675
rect 1903 4641 1912 4675
rect 1860 4632 1912 4641
rect 2504 4632 2556 4684
rect 3240 4564 3292 4616
rect 3424 4564 3476 4616
rect 4436 4700 4488 4752
rect 4712 4632 4764 4684
rect 4068 4428 4120 4480
rect 4160 4428 4212 4480
rect 4620 4564 4672 4616
rect 4988 4564 5040 4616
rect 6276 4632 6328 4684
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 6092 4564 6144 4573
rect 7840 4564 7892 4616
rect 8300 4564 8352 4616
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 12808 4768 12860 4820
rect 13912 4768 13964 4820
rect 14280 4768 14332 4820
rect 14372 4768 14424 4820
rect 8944 4675 8996 4684
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 9220 4675 9272 4684
rect 9220 4641 9229 4675
rect 9229 4641 9263 4675
rect 9263 4641 9272 4675
rect 9220 4632 9272 4641
rect 11520 4700 11572 4752
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 10784 4607 10836 4616
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 10784 4564 10836 4573
rect 11152 4607 11204 4616
rect 11152 4573 11161 4607
rect 11161 4573 11195 4607
rect 11195 4573 11204 4607
rect 11152 4564 11204 4573
rect 11520 4607 11572 4616
rect 11520 4573 11529 4607
rect 11529 4573 11563 4607
rect 11563 4573 11572 4607
rect 11520 4564 11572 4573
rect 5540 4471 5592 4480
rect 5540 4437 5549 4471
rect 5549 4437 5583 4471
rect 5583 4437 5592 4471
rect 5540 4428 5592 4437
rect 8300 4471 8352 4480
rect 8300 4437 8309 4471
rect 8309 4437 8343 4471
rect 8343 4437 8352 4471
rect 8300 4428 8352 4437
rect 8576 4471 8628 4480
rect 8576 4437 8585 4471
rect 8585 4437 8619 4471
rect 8619 4437 8628 4471
rect 8576 4428 8628 4437
rect 10508 4496 10560 4548
rect 10692 4496 10744 4548
rect 12624 4564 12676 4616
rect 14004 4564 14056 4616
rect 14096 4496 14148 4548
rect 15016 4607 15068 4616
rect 15016 4573 15025 4607
rect 15025 4573 15059 4607
rect 15059 4573 15068 4607
rect 15016 4564 15068 4573
rect 15108 4564 15160 4616
rect 15476 4496 15528 4548
rect 11336 4428 11388 4480
rect 11428 4428 11480 4480
rect 11612 4471 11664 4480
rect 11612 4437 11621 4471
rect 11621 4437 11655 4471
rect 11655 4437 11664 4471
rect 11612 4428 11664 4437
rect 12440 4428 12492 4480
rect 12716 4471 12768 4480
rect 12716 4437 12725 4471
rect 12725 4437 12759 4471
rect 12759 4437 12768 4471
rect 12716 4428 12768 4437
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 13728 4471 13780 4480
rect 13728 4437 13737 4471
rect 13737 4437 13771 4471
rect 13771 4437 13780 4471
rect 13728 4428 13780 4437
rect 14188 4428 14240 4480
rect 15660 4471 15712 4480
rect 15660 4437 15669 4471
rect 15669 4437 15703 4471
rect 15703 4437 15712 4471
rect 15660 4428 15712 4437
rect 3473 4326 3525 4378
rect 3537 4326 3589 4378
rect 3601 4326 3653 4378
rect 3665 4326 3717 4378
rect 3729 4326 3781 4378
rect 7199 4326 7251 4378
rect 7263 4326 7315 4378
rect 7327 4326 7379 4378
rect 7391 4326 7443 4378
rect 7455 4326 7507 4378
rect 10925 4326 10977 4378
rect 10989 4326 11041 4378
rect 11053 4326 11105 4378
rect 11117 4326 11169 4378
rect 11181 4326 11233 4378
rect 14651 4326 14703 4378
rect 14715 4326 14767 4378
rect 14779 4326 14831 4378
rect 14843 4326 14895 4378
rect 14907 4326 14959 4378
rect 3884 4224 3936 4276
rect 4068 4267 4120 4276
rect 4068 4233 4077 4267
rect 4077 4233 4111 4267
rect 4111 4233 4120 4267
rect 4068 4224 4120 4233
rect 4436 4224 4488 4276
rect 5448 4224 5500 4276
rect 6092 4224 6144 4276
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 3240 4088 3292 4140
rect 3792 4156 3844 4208
rect 3148 4020 3200 4072
rect 3332 4020 3384 4072
rect 4068 4088 4120 4140
rect 4620 4156 4672 4208
rect 9128 4224 9180 4276
rect 11428 4224 11480 4276
rect 6276 4088 6328 4140
rect 7748 4088 7800 4140
rect 8300 4088 8352 4140
rect 8944 4088 8996 4140
rect 9496 4131 9548 4140
rect 9496 4097 9505 4131
rect 9505 4097 9539 4131
rect 9539 4097 9548 4131
rect 9496 4088 9548 4097
rect 3332 3884 3384 3936
rect 4528 4063 4580 4072
rect 4528 4029 4537 4063
rect 4537 4029 4571 4063
rect 4571 4029 4580 4063
rect 4528 4020 4580 4029
rect 6092 3884 6144 3936
rect 8576 4020 8628 4072
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 10508 4020 10560 4072
rect 11336 4088 11388 4140
rect 14188 4224 14240 4276
rect 14280 4224 14332 4276
rect 15016 4224 15068 4276
rect 15476 4267 15528 4276
rect 15476 4233 15485 4267
rect 15485 4233 15519 4267
rect 15519 4233 15528 4267
rect 15476 4224 15528 4233
rect 12716 4156 12768 4208
rect 13912 4156 13964 4208
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 11704 4020 11756 4072
rect 12440 4020 12492 4072
rect 12624 4131 12676 4140
rect 12624 4097 12633 4131
rect 12633 4097 12667 4131
rect 12667 4097 12676 4131
rect 12624 4088 12676 4097
rect 12808 4088 12860 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 14556 4088 14608 4140
rect 13728 4020 13780 4072
rect 14464 4020 14516 4072
rect 14924 4020 14976 4072
rect 15292 4063 15344 4072
rect 15292 4029 15301 4063
rect 15301 4029 15335 4063
rect 15335 4029 15344 4063
rect 15292 4020 15344 4029
rect 11336 3952 11388 4004
rect 12164 3952 12216 4004
rect 12716 3952 12768 4004
rect 6460 3884 6512 3936
rect 8300 3884 8352 3936
rect 2813 3782 2865 3834
rect 2877 3782 2929 3834
rect 2941 3782 2993 3834
rect 3005 3782 3057 3834
rect 3069 3782 3121 3834
rect 6539 3782 6591 3834
rect 6603 3782 6655 3834
rect 6667 3782 6719 3834
rect 6731 3782 6783 3834
rect 6795 3782 6847 3834
rect 10265 3782 10317 3834
rect 10329 3782 10381 3834
rect 10393 3782 10445 3834
rect 10457 3782 10509 3834
rect 10521 3782 10573 3834
rect 13991 3782 14043 3834
rect 14055 3782 14107 3834
rect 14119 3782 14171 3834
rect 14183 3782 14235 3834
rect 14247 3782 14299 3834
rect 4528 3680 4580 3732
rect 5540 3680 5592 3732
rect 6092 3723 6144 3732
rect 6092 3689 6101 3723
rect 6101 3689 6135 3723
rect 6135 3689 6144 3723
rect 6092 3680 6144 3689
rect 6276 3680 6328 3732
rect 7656 3680 7708 3732
rect 7932 3723 7984 3732
rect 7932 3689 7941 3723
rect 7941 3689 7975 3723
rect 7975 3689 7984 3723
rect 7932 3680 7984 3689
rect 9864 3680 9916 3732
rect 9956 3680 10008 3732
rect 11704 3680 11756 3732
rect 13636 3680 13688 3732
rect 13912 3723 13964 3732
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 14924 3680 14976 3732
rect 15292 3680 15344 3732
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 4988 3612 5040 3664
rect 3240 3476 3292 3528
rect 2136 3451 2188 3460
rect 2136 3417 2145 3451
rect 2145 3417 2179 3451
rect 2179 3417 2188 3451
rect 2136 3408 2188 3417
rect 3884 3340 3936 3392
rect 5448 3476 5500 3528
rect 11520 3612 11572 3664
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 7748 3476 7800 3528
rect 7932 3476 7984 3528
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 9496 3544 9548 3596
rect 12992 3544 13044 3596
rect 5172 3340 5224 3392
rect 11336 3476 11388 3528
rect 11980 3519 12032 3528
rect 10600 3340 10652 3392
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 14004 3476 14056 3528
rect 15108 3476 15160 3528
rect 15016 3408 15068 3460
rect 3473 3238 3525 3290
rect 3537 3238 3589 3290
rect 3601 3238 3653 3290
rect 3665 3238 3717 3290
rect 3729 3238 3781 3290
rect 7199 3238 7251 3290
rect 7263 3238 7315 3290
rect 7327 3238 7379 3290
rect 7391 3238 7443 3290
rect 7455 3238 7507 3290
rect 10925 3238 10977 3290
rect 10989 3238 11041 3290
rect 11053 3238 11105 3290
rect 11117 3238 11169 3290
rect 11181 3238 11233 3290
rect 14651 3238 14703 3290
rect 14715 3238 14767 3290
rect 14779 3238 14831 3290
rect 14843 3238 14895 3290
rect 14907 3238 14959 3290
rect 2136 3136 2188 3188
rect 3884 3136 3936 3188
rect 5632 3136 5684 3188
rect 7932 3136 7984 3188
rect 9772 3136 9824 3188
rect 10784 3136 10836 3188
rect 11980 3136 12032 3188
rect 12072 3136 12124 3188
rect 12624 3136 12676 3188
rect 12808 3136 12860 3188
rect 2780 3000 2832 3052
rect 3332 3068 3384 3120
rect 5908 3068 5960 3120
rect 6460 3000 6512 3052
rect 1676 2932 1728 2984
rect 7104 3000 7156 3052
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 8300 2864 8352 2916
rect 4436 2796 4488 2848
rect 11428 3000 11480 3052
rect 11612 3000 11664 3052
rect 14372 3136 14424 3188
rect 15016 3136 15068 3188
rect 14004 3068 14056 3120
rect 12992 3000 13044 3052
rect 10600 2864 10652 2916
rect 13912 2932 13964 2984
rect 14556 2932 14608 2984
rect 15660 3000 15712 3052
rect 14740 2864 14792 2916
rect 12072 2796 12124 2848
rect 12440 2796 12492 2848
rect 15108 2796 15160 2848
rect 2813 2694 2865 2746
rect 2877 2694 2929 2746
rect 2941 2694 2993 2746
rect 3005 2694 3057 2746
rect 3069 2694 3121 2746
rect 6539 2694 6591 2746
rect 6603 2694 6655 2746
rect 6667 2694 6719 2746
rect 6731 2694 6783 2746
rect 6795 2694 6847 2746
rect 10265 2694 10317 2746
rect 10329 2694 10381 2746
rect 10393 2694 10445 2746
rect 10457 2694 10509 2746
rect 10521 2694 10573 2746
rect 13991 2694 14043 2746
rect 14055 2694 14107 2746
rect 14119 2694 14171 2746
rect 14183 2694 14235 2746
rect 14247 2694 14299 2746
rect 13176 2592 13228 2644
rect 1676 2567 1728 2576
rect 1676 2533 1685 2567
rect 1685 2533 1719 2567
rect 1719 2533 1728 2567
rect 1676 2524 1728 2533
rect 14740 2567 14792 2576
rect 14740 2533 14749 2567
rect 14749 2533 14783 2567
rect 14783 2533 14792 2567
rect 14740 2524 14792 2533
rect 15108 2499 15160 2508
rect 15108 2465 15117 2499
rect 15117 2465 15151 2499
rect 15151 2465 15160 2499
rect 15108 2456 15160 2465
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 12716 2388 12768 2440
rect 20 2320 72 2372
rect 9680 2252 9732 2304
rect 12900 2252 12952 2304
rect 3473 2150 3525 2202
rect 3537 2150 3589 2202
rect 3601 2150 3653 2202
rect 3665 2150 3717 2202
rect 3729 2150 3781 2202
rect 7199 2150 7251 2202
rect 7263 2150 7315 2202
rect 7327 2150 7379 2202
rect 7391 2150 7443 2202
rect 7455 2150 7507 2202
rect 10925 2150 10977 2202
rect 10989 2150 11041 2202
rect 11053 2150 11105 2202
rect 11117 2150 11169 2202
rect 11181 2150 11233 2202
rect 14651 2150 14703 2202
rect 14715 2150 14767 2202
rect 14779 2150 14831 2202
rect 14843 2150 14895 2202
rect 14907 2150 14959 2202
<< metal2 >>
rect 662 18546 718 19346
rect 3882 18546 3938 19346
rect 7102 18546 7158 19346
rect 10322 18546 10378 19346
rect 13542 18546 13598 19346
rect 16762 18546 16818 19346
rect 676 9625 704 18546
rect 2813 16892 3121 16901
rect 2813 16890 2819 16892
rect 2875 16890 2899 16892
rect 2955 16890 2979 16892
rect 3035 16890 3059 16892
rect 3115 16890 3121 16892
rect 2875 16838 2877 16890
rect 3057 16838 3059 16890
rect 2813 16836 2819 16838
rect 2875 16836 2899 16838
rect 2955 16836 2979 16838
rect 3035 16836 3059 16838
rect 3115 16836 3121 16838
rect 2813 16827 3121 16836
rect 6539 16892 6847 16901
rect 6539 16890 6545 16892
rect 6601 16890 6625 16892
rect 6681 16890 6705 16892
rect 6761 16890 6785 16892
rect 6841 16890 6847 16892
rect 6601 16838 6603 16890
rect 6783 16838 6785 16890
rect 6539 16836 6545 16838
rect 6601 16836 6625 16838
rect 6681 16836 6705 16838
rect 6761 16836 6785 16838
rect 6841 16836 6847 16838
rect 6539 16827 6847 16836
rect 10265 16892 10573 16901
rect 10265 16890 10271 16892
rect 10327 16890 10351 16892
rect 10407 16890 10431 16892
rect 10487 16890 10511 16892
rect 10567 16890 10573 16892
rect 10327 16838 10329 16890
rect 10509 16838 10511 16890
rect 10265 16836 10271 16838
rect 10327 16836 10351 16838
rect 10407 16836 10431 16838
rect 10487 16836 10511 16838
rect 10567 16836 10573 16838
rect 10265 16827 10573 16836
rect 13991 16892 14299 16901
rect 13991 16890 13997 16892
rect 14053 16890 14077 16892
rect 14133 16890 14157 16892
rect 14213 16890 14237 16892
rect 14293 16890 14299 16892
rect 14053 16838 14055 16890
rect 14235 16838 14237 16890
rect 13991 16836 13997 16838
rect 14053 16836 14077 16838
rect 14133 16836 14157 16838
rect 14213 16836 14237 16838
rect 14293 16836 14299 16838
rect 13991 16827 14299 16836
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 4344 16448 4396 16454
rect 4344 16390 4396 16396
rect 3473 16348 3781 16357
rect 3473 16346 3479 16348
rect 3535 16346 3559 16348
rect 3615 16346 3639 16348
rect 3695 16346 3719 16348
rect 3775 16346 3781 16348
rect 3535 16294 3537 16346
rect 3717 16294 3719 16346
rect 3473 16292 3479 16294
rect 3535 16292 3559 16294
rect 3615 16292 3639 16294
rect 3695 16292 3719 16294
rect 3775 16292 3781 16294
rect 3473 16283 3781 16292
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 2813 15804 3121 15813
rect 2813 15802 2819 15804
rect 2875 15802 2899 15804
rect 2955 15802 2979 15804
rect 3035 15802 3059 15804
rect 3115 15802 3121 15804
rect 2875 15750 2877 15802
rect 3057 15750 3059 15802
rect 2813 15748 2819 15750
rect 2875 15748 2899 15750
rect 2955 15748 2979 15750
rect 3035 15748 3059 15750
rect 3115 15748 3121 15750
rect 2813 15739 3121 15748
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2792 14890 2820 15302
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2700 13938 2728 14758
rect 2813 14716 3121 14725
rect 2813 14714 2819 14716
rect 2875 14714 2899 14716
rect 2955 14714 2979 14716
rect 3035 14714 3059 14716
rect 3115 14714 3121 14716
rect 2875 14662 2877 14714
rect 3057 14662 3059 14714
rect 2813 14660 2819 14662
rect 2875 14660 2899 14662
rect 2955 14660 2979 14662
rect 3035 14660 3059 14662
rect 3115 14660 3121 14662
rect 2813 14651 3121 14660
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2516 13394 2544 13670
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1964 12646 1992 13126
rect 2700 12782 2728 13874
rect 2813 13628 3121 13637
rect 2813 13626 2819 13628
rect 2875 13626 2899 13628
rect 2955 13626 2979 13628
rect 3035 13626 3059 13628
rect 3115 13626 3121 13628
rect 2875 13574 2877 13626
rect 3057 13574 3059 13626
rect 2813 13572 2819 13574
rect 2875 13572 2899 13574
rect 2955 13572 2979 13574
rect 3035 13572 3059 13574
rect 3115 13572 3121 13574
rect 2813 13563 3121 13572
rect 3160 13326 3188 15370
rect 3473 15260 3781 15269
rect 3473 15258 3479 15260
rect 3535 15258 3559 15260
rect 3615 15258 3639 15260
rect 3695 15258 3719 15260
rect 3775 15258 3781 15260
rect 3535 15206 3537 15258
rect 3717 15206 3719 15258
rect 3473 15204 3479 15206
rect 3535 15204 3559 15206
rect 3615 15204 3639 15206
rect 3695 15204 3719 15206
rect 3775 15204 3781 15206
rect 3473 15195 3781 15204
rect 3896 15162 3924 15982
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 4264 15026 4292 15302
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 3988 14906 4016 14962
rect 4356 14958 4384 16390
rect 5368 16250 5396 16526
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7116 16250 7144 16390
rect 7199 16348 7507 16357
rect 7199 16346 7205 16348
rect 7261 16346 7285 16348
rect 7341 16346 7365 16348
rect 7421 16346 7445 16348
rect 7501 16346 7507 16348
rect 7261 16294 7263 16346
rect 7443 16294 7445 16346
rect 7199 16292 7205 16294
rect 7261 16292 7285 16294
rect 7341 16292 7365 16294
rect 7421 16292 7445 16294
rect 7501 16292 7507 16294
rect 7199 16283 7507 16292
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4632 15570 4660 15846
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4632 15094 4660 15506
rect 5000 15094 5028 16186
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5080 15904 5132 15910
rect 5080 15846 5132 15852
rect 5092 15706 5120 15846
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 4344 14952 4396 14958
rect 3988 14878 4200 14906
rect 4344 14894 4396 14900
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 3473 14172 3781 14181
rect 3473 14170 3479 14172
rect 3535 14170 3559 14172
rect 3615 14170 3639 14172
rect 3695 14170 3719 14172
rect 3775 14170 3781 14172
rect 3535 14118 3537 14170
rect 3717 14118 3719 14170
rect 3473 14116 3479 14118
rect 3535 14116 3559 14118
rect 3615 14116 3639 14118
rect 3695 14116 3719 14118
rect 3775 14116 3781 14118
rect 3473 14107 3781 14116
rect 4172 14074 4200 14878
rect 4724 14618 4752 14894
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 12102 1992 12582
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1964 11626 1992 12038
rect 2148 11898 2176 12718
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2700 11762 2728 12718
rect 2884 12646 2912 12854
rect 3068 12730 3096 13126
rect 3160 12986 3188 13262
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3068 12702 3280 12730
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 2813 12540 3121 12549
rect 2813 12538 2819 12540
rect 2875 12538 2899 12540
rect 2955 12538 2979 12540
rect 3035 12538 3059 12540
rect 3115 12538 3121 12540
rect 2875 12486 2877 12538
rect 3057 12486 3059 12538
rect 2813 12484 2819 12486
rect 2875 12484 2899 12486
rect 2955 12484 2979 12486
rect 3035 12484 3059 12486
rect 3115 12484 3121 12486
rect 2813 12475 3121 12484
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 3160 11642 3188 12582
rect 3252 11830 3280 12702
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 3344 11762 3372 13262
rect 3896 13190 3924 13806
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3473 13084 3781 13093
rect 3473 13082 3479 13084
rect 3535 13082 3559 13084
rect 3615 13082 3639 13084
rect 3695 13082 3719 13084
rect 3775 13082 3781 13084
rect 3535 13030 3537 13082
rect 3717 13030 3719 13082
rect 3473 13028 3479 13030
rect 3535 13028 3559 13030
rect 3615 13028 3639 13030
rect 3695 13028 3719 13030
rect 3775 13028 3781 13030
rect 3473 13019 3781 13028
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3436 12170 3464 12922
rect 3896 12714 3924 13126
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3473 11996 3781 12005
rect 3473 11994 3479 11996
rect 3535 11994 3559 11996
rect 3615 11994 3639 11996
rect 3695 11994 3719 11996
rect 3775 11994 3781 11996
rect 3535 11942 3537 11994
rect 3717 11942 3719 11994
rect 3473 11940 3479 11942
rect 3535 11940 3559 11942
rect 3615 11940 3639 11942
rect 3695 11940 3719 11942
rect 3775 11940 3781 11942
rect 3473 11931 3781 11940
rect 3896 11898 3924 12242
rect 3976 12164 4028 12170
rect 3976 12106 4028 12112
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3988 11830 4016 12106
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 2700 11614 3188 11642
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10305 980 10610
rect 1964 10606 1992 11562
rect 2700 11268 2728 11614
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 2813 11452 3121 11461
rect 2813 11450 2819 11452
rect 2875 11450 2899 11452
rect 2955 11450 2979 11452
rect 3035 11450 3059 11452
rect 3115 11450 3121 11452
rect 2875 11398 2877 11450
rect 3057 11398 3059 11450
rect 2813 11396 2819 11398
rect 2875 11396 2899 11398
rect 2955 11396 2979 11398
rect 3035 11396 3059 11398
rect 3115 11396 3121 11398
rect 2813 11387 3121 11396
rect 2700 11240 2912 11268
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 2228 10600 2280 10606
rect 2792 10554 2820 10950
rect 2884 10742 2912 11240
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2976 10606 3004 10950
rect 3160 10810 3188 11494
rect 3252 11286 3280 11630
rect 3528 11626 3556 11766
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3792 11620 3844 11626
rect 3792 11562 3844 11568
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 2228 10542 2280 10548
rect 938 10296 994 10305
rect 2240 10266 2268 10542
rect 2700 10526 2820 10554
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 938 10231 994 10240
rect 2228 10260 2280 10266
rect 2700 10248 2728 10526
rect 2813 10364 3121 10373
rect 2813 10362 2819 10364
rect 2875 10362 2899 10364
rect 2955 10362 2979 10364
rect 3035 10362 3059 10364
rect 3115 10362 3121 10364
rect 2875 10310 2877 10362
rect 3057 10310 3059 10362
rect 2813 10308 2819 10310
rect 2875 10308 2899 10310
rect 2955 10308 2979 10310
rect 3035 10308 3059 10310
rect 3115 10308 3121 10310
rect 2813 10299 3121 10308
rect 2700 10220 2820 10248
rect 2228 10202 2280 10208
rect 2792 10062 2820 10220
rect 3160 10130 3188 10746
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 3252 9926 3280 11018
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3344 9704 3372 11290
rect 3804 10962 3832 11562
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3896 11132 3924 11494
rect 3988 11286 4016 11766
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4080 11226 4108 11494
rect 4172 11354 4200 14010
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4356 12850 4384 13262
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4356 11694 4384 12786
rect 4632 12102 4660 13874
rect 4816 12850 4844 14010
rect 5000 14006 5028 15030
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5276 14414 5304 14758
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5460 14074 5488 14758
rect 5552 14550 5580 15982
rect 6012 15502 6040 16050
rect 6539 15804 6847 15813
rect 6539 15802 6545 15804
rect 6601 15802 6625 15804
rect 6681 15802 6705 15804
rect 6761 15802 6785 15804
rect 6841 15802 6847 15804
rect 6601 15750 6603 15802
rect 6783 15750 6785 15802
rect 6539 15748 6545 15750
rect 6601 15748 6625 15750
rect 6681 15748 6705 15750
rect 6761 15748 6785 15750
rect 6841 15748 6847 15750
rect 6539 15739 6847 15748
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5540 14408 5592 14414
rect 5644 14396 5672 15302
rect 6012 15026 6040 15438
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6380 15162 6408 15302
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6564 15026 6592 15302
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 5592 14368 5672 14396
rect 5540 14350 5592 14356
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 4988 14000 5040 14006
rect 4988 13942 5040 13948
rect 5552 13938 5580 14350
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5736 14074 5764 14214
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 5000 12434 5028 12922
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 4816 12406 5028 12434
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4264 11354 4292 11630
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 11354 4384 11494
rect 4448 11354 4476 11698
rect 4540 11354 4568 12038
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4068 11220 4120 11226
rect 4068 11162 4120 11168
rect 4344 11144 4396 11150
rect 3896 11104 4344 11132
rect 4632 11132 4660 12038
rect 4724 11694 4752 12038
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4816 11218 4844 12406
rect 5092 12102 5120 12786
rect 5184 12730 5212 12786
rect 5184 12702 5304 12730
rect 5276 12434 5304 12702
rect 5460 12434 5488 12786
rect 5920 12782 5948 14214
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6012 12714 6040 14962
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6196 14550 6224 14758
rect 6539 14716 6847 14725
rect 6539 14714 6545 14716
rect 6601 14714 6625 14716
rect 6681 14714 6705 14716
rect 6761 14714 6785 14716
rect 6841 14714 6847 14716
rect 6601 14662 6603 14714
rect 6783 14662 6785 14714
rect 6539 14660 6545 14662
rect 6601 14660 6625 14662
rect 6681 14660 6705 14662
rect 6761 14660 6785 14662
rect 6841 14660 6847 14662
rect 6539 14651 6847 14660
rect 6184 14544 6236 14550
rect 6184 14486 6236 14492
rect 6539 13628 6847 13637
rect 6539 13626 6545 13628
rect 6601 13626 6625 13628
rect 6681 13626 6705 13628
rect 6761 13626 6785 13628
rect 6841 13626 6847 13628
rect 6601 13574 6603 13626
rect 6783 13574 6785 13626
rect 6539 13572 6545 13574
rect 6601 13572 6625 13574
rect 6681 13572 6705 13574
rect 6761 13572 6785 13574
rect 6841 13572 6847 13574
rect 6539 13563 6847 13572
rect 6932 13326 6960 15438
rect 7199 15260 7507 15269
rect 7199 15258 7205 15260
rect 7261 15258 7285 15260
rect 7341 15258 7365 15260
rect 7421 15258 7445 15260
rect 7501 15258 7507 15260
rect 7261 15206 7263 15258
rect 7443 15206 7445 15258
rect 7199 15204 7205 15206
rect 7261 15204 7285 15206
rect 7341 15204 7365 15206
rect 7421 15204 7445 15206
rect 7501 15204 7507 15206
rect 7199 15195 7507 15204
rect 7668 15162 7696 16526
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7852 15706 7880 15846
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7944 15570 7972 15982
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7380 15088 7432 15094
rect 7380 15030 7432 15036
rect 8128 15042 8156 16594
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8220 15706 8248 15982
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8404 15162 8432 16594
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 9140 16250 9168 16390
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8496 15162 8524 15438
rect 9140 15162 9168 16186
rect 10796 16182 10824 16390
rect 10925 16348 11233 16357
rect 10925 16346 10931 16348
rect 10987 16346 11011 16348
rect 11067 16346 11091 16348
rect 11147 16346 11171 16348
rect 11227 16346 11233 16348
rect 10987 16294 10989 16346
rect 11169 16294 11171 16346
rect 10925 16292 10931 16294
rect 10987 16292 11011 16294
rect 11067 16292 11091 16294
rect 11147 16292 11171 16294
rect 11227 16292 11233 16294
rect 10925 16283 11233 16292
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10152 15706 10180 16118
rect 10265 15804 10573 15813
rect 10265 15802 10271 15804
rect 10327 15802 10351 15804
rect 10407 15802 10431 15804
rect 10487 15802 10511 15804
rect 10567 15802 10573 15804
rect 10327 15750 10329 15802
rect 10509 15750 10511 15802
rect 10265 15748 10271 15750
rect 10327 15748 10351 15750
rect 10407 15748 10431 15750
rect 10487 15748 10511 15750
rect 10567 15748 10573 15750
rect 10265 15739 10573 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14618 7328 14758
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7392 14550 7420 15030
rect 8128 15026 8432 15042
rect 8128 15020 8444 15026
rect 8128 15014 8392 15020
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7484 14618 7512 14894
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7392 14414 7420 14486
rect 8220 14414 8248 15014
rect 8392 14962 8444 14968
rect 9140 14618 9168 15098
rect 9692 15094 9720 15302
rect 9784 15094 9812 15438
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9508 14482 9536 14758
rect 9784 14482 9812 15030
rect 9876 14618 9904 15438
rect 10152 15094 10180 15642
rect 11348 15502 11376 16526
rect 11440 16250 11468 16594
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 12360 16046 12388 16526
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15570 12204 15846
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 10925 15260 11233 15269
rect 10925 15258 10931 15260
rect 10987 15258 11011 15260
rect 11067 15258 11091 15260
rect 11147 15258 11171 15260
rect 11227 15258 11233 15260
rect 10987 15206 10989 15258
rect 11169 15206 11171 15258
rect 10925 15204 10931 15206
rect 10987 15204 11011 15206
rect 11067 15204 11091 15206
rect 11147 15204 11171 15206
rect 11227 15204 11233 15206
rect 10925 15195 11233 15204
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5184 12406 5304 12434
rect 5368 12406 5488 12434
rect 5184 12238 5212 12406
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 5092 11150 5120 12038
rect 4712 11144 4764 11150
rect 4632 11104 4712 11132
rect 4344 11086 4396 11092
rect 4712 11086 4764 11092
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4252 11008 4304 11014
rect 3804 10934 4016 10962
rect 5184 10996 5212 12174
rect 5276 11354 5304 12174
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5368 11014 5396 12406
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 11200 5488 11630
rect 5552 11354 5580 12582
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 6012 11218 6040 12650
rect 6472 12434 6500 12718
rect 6539 12540 6847 12549
rect 6539 12538 6545 12540
rect 6601 12538 6625 12540
rect 6681 12538 6705 12540
rect 6761 12538 6785 12540
rect 6841 12538 6847 12540
rect 6601 12486 6603 12538
rect 6783 12486 6785 12538
rect 6539 12484 6545 12486
rect 6601 12484 6625 12486
rect 6681 12484 6705 12486
rect 6761 12484 6785 12486
rect 6841 12484 6847 12486
rect 6539 12475 6847 12484
rect 6552 12436 6604 12442
rect 6472 12406 6552 12434
rect 6932 12434 6960 13262
rect 6552 12378 6604 12384
rect 6840 12406 6960 12434
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6196 11898 6224 12174
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6748 11694 6776 12038
rect 6840 11830 6868 12406
rect 7024 12374 7052 14214
rect 7199 14172 7507 14181
rect 7199 14170 7205 14172
rect 7261 14170 7285 14172
rect 7341 14170 7365 14172
rect 7421 14170 7445 14172
rect 7501 14170 7507 14172
rect 7261 14118 7263 14170
rect 7443 14118 7445 14170
rect 7199 14116 7205 14118
rect 7261 14116 7285 14118
rect 7341 14116 7365 14118
rect 7421 14116 7445 14118
rect 7501 14116 7507 14118
rect 7199 14107 7507 14116
rect 7944 14074 7972 14214
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 8300 13252 8352 13258
rect 8300 13194 8352 13200
rect 7199 13084 7507 13093
rect 7199 13082 7205 13084
rect 7261 13082 7285 13084
rect 7341 13082 7365 13084
rect 7421 13082 7445 13084
rect 7501 13082 7507 13084
rect 7261 13030 7263 13082
rect 7443 13030 7445 13082
rect 7199 13028 7205 13030
rect 7261 13028 7285 13030
rect 7341 13028 7365 13030
rect 7421 13028 7445 13030
rect 7501 13028 7507 13030
rect 7199 13019 7507 13028
rect 7576 12986 7604 13194
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6539 11452 6847 11461
rect 6539 11450 6545 11452
rect 6601 11450 6625 11452
rect 6681 11450 6705 11452
rect 6761 11450 6785 11452
rect 6841 11450 6847 11452
rect 6601 11398 6603 11450
rect 6783 11398 6785 11450
rect 6539 11396 6545 11398
rect 6601 11396 6625 11398
rect 6681 11396 6705 11398
rect 6761 11396 6785 11398
rect 6841 11396 6847 11398
rect 6539 11387 6847 11396
rect 7024 11286 7052 12310
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 5540 11212 5592 11218
rect 5460 11172 5540 11200
rect 5540 11154 5592 11160
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 4252 10950 4304 10956
rect 5000 10968 5212 10996
rect 5356 11008 5408 11014
rect 3473 10908 3781 10917
rect 3473 10906 3479 10908
rect 3535 10906 3559 10908
rect 3615 10906 3639 10908
rect 3695 10906 3719 10908
rect 3775 10906 3781 10908
rect 3535 10854 3537 10906
rect 3717 10854 3719 10906
rect 3473 10852 3479 10854
rect 3535 10852 3559 10854
rect 3615 10852 3639 10854
rect 3695 10852 3719 10854
rect 3775 10852 3781 10854
rect 3473 10843 3781 10852
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3804 10266 3832 10406
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3473 9820 3781 9829
rect 3473 9818 3479 9820
rect 3535 9818 3559 9820
rect 3615 9818 3639 9820
rect 3695 9818 3719 9820
rect 3775 9818 3781 9820
rect 3535 9766 3537 9818
rect 3717 9766 3719 9818
rect 3473 9764 3479 9766
rect 3535 9764 3559 9766
rect 3615 9764 3639 9766
rect 3695 9764 3719 9766
rect 3775 9764 3781 9766
rect 3473 9755 3781 9764
rect 3896 9738 3924 9998
rect 3252 9676 3372 9704
rect 3804 9710 3924 9738
rect 3148 9648 3200 9654
rect 662 9616 718 9625
rect 3148 9590 3200 9596
rect 662 9551 718 9560
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1872 8498 1900 8910
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 7410 1900 8434
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1872 6866 1900 7346
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 1872 4690 1900 6802
rect 2700 5710 2728 9318
rect 2813 9276 3121 9285
rect 2813 9274 2819 9276
rect 2875 9274 2899 9276
rect 2955 9274 2979 9276
rect 3035 9274 3059 9276
rect 3115 9274 3121 9276
rect 2875 9222 2877 9274
rect 3057 9222 3059 9274
rect 2813 9220 2819 9222
rect 2875 9220 2899 9222
rect 2955 9220 2979 9222
rect 3035 9220 3059 9222
rect 3115 9220 3121 9222
rect 2813 9211 3121 9220
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 8566 3096 8774
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2813 8188 3121 8197
rect 2813 8186 2819 8188
rect 2875 8186 2899 8188
rect 2955 8186 2979 8188
rect 3035 8186 3059 8188
rect 3115 8186 3121 8188
rect 2875 8134 2877 8186
rect 3057 8134 3059 8186
rect 2813 8132 2819 8134
rect 2875 8132 2899 8134
rect 2955 8132 2979 8134
rect 3035 8132 3059 8134
rect 3115 8132 3121 8134
rect 2813 8123 3121 8132
rect 2813 7100 3121 7109
rect 2813 7098 2819 7100
rect 2875 7098 2899 7100
rect 2955 7098 2979 7100
rect 3035 7098 3059 7100
rect 3115 7098 3121 7100
rect 2875 7046 2877 7098
rect 3057 7046 3059 7098
rect 2813 7044 2819 7046
rect 2875 7044 2899 7046
rect 2955 7044 2979 7046
rect 3035 7044 3059 7046
rect 3115 7044 3121 7046
rect 2813 7035 3121 7044
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6202 3096 6598
rect 3160 6322 3188 9590
rect 3252 8974 3280 9676
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8294 3280 8910
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3252 7546 3280 8230
rect 3344 7886 3372 9522
rect 3804 9382 3832 9710
rect 3988 9586 4016 10934
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 4080 9586 4108 9930
rect 4172 9926 4200 10610
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4172 9722 4200 9862
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3473 8732 3781 8741
rect 3473 8730 3479 8732
rect 3535 8730 3559 8732
rect 3615 8730 3639 8732
rect 3695 8730 3719 8732
rect 3775 8730 3781 8732
rect 3535 8678 3537 8730
rect 3717 8678 3719 8730
rect 3473 8676 3479 8678
rect 3535 8676 3559 8678
rect 3615 8676 3639 8678
rect 3695 8676 3719 8678
rect 3775 8676 3781 8678
rect 3473 8667 3781 8676
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3252 6798 3280 7482
rect 3344 7188 3372 7686
rect 3473 7644 3781 7653
rect 3473 7642 3479 7644
rect 3535 7642 3559 7644
rect 3615 7642 3639 7644
rect 3695 7642 3719 7644
rect 3775 7642 3781 7644
rect 3535 7590 3537 7642
rect 3717 7590 3719 7642
rect 3473 7588 3479 7590
rect 3535 7588 3559 7590
rect 3615 7588 3639 7590
rect 3695 7588 3719 7590
rect 3775 7588 3781 7590
rect 3473 7579 3781 7588
rect 3896 7410 3924 9522
rect 4080 9466 4108 9522
rect 3988 9438 4108 9466
rect 3988 8090 4016 9438
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 9178 4108 9318
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3424 7200 3476 7206
rect 3344 7160 3424 7188
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3068 6174 3188 6202
rect 2813 6012 3121 6021
rect 2813 6010 2819 6012
rect 2875 6010 2899 6012
rect 2955 6010 2979 6012
rect 3035 6010 3059 6012
rect 3115 6010 3121 6012
rect 2875 5958 2877 6010
rect 3057 5958 3059 6010
rect 2813 5956 2819 5958
rect 2875 5956 2899 5958
rect 2955 5956 2979 5958
rect 3035 5956 3059 5958
rect 3115 5956 3121 5958
rect 2813 5947 3121 5956
rect 3160 5828 3188 6174
rect 3068 5800 3188 5828
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 2792 5114 2820 5578
rect 3068 5234 3096 5800
rect 3252 5710 3280 6326
rect 3344 6322 3372 7160
rect 3424 7142 3476 7148
rect 3988 6746 4016 7686
rect 4080 6934 4108 7822
rect 4172 7342 4200 9658
rect 4264 7546 4292 10950
rect 5000 10674 5028 10968
rect 5356 10950 5408 10956
rect 5368 10674 5396 10950
rect 5552 10674 5580 11154
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4632 9518 4660 10542
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 9586 5212 10406
rect 5552 10266 5580 10610
rect 6539 10364 6847 10373
rect 6539 10362 6545 10364
rect 6601 10362 6625 10364
rect 6681 10362 6705 10364
rect 6761 10362 6785 10364
rect 6841 10362 6847 10364
rect 6601 10310 6603 10362
rect 6783 10310 6785 10362
rect 6539 10308 6545 10310
rect 6601 10308 6625 10310
rect 6681 10308 6705 10310
rect 6761 10308 6785 10310
rect 6841 10308 6847 10310
rect 6539 10299 6847 10308
rect 7116 10266 7144 12786
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7199 11996 7507 12005
rect 7199 11994 7205 11996
rect 7261 11994 7285 11996
rect 7341 11994 7365 11996
rect 7421 11994 7445 11996
rect 7501 11994 7507 11996
rect 7261 11942 7263 11994
rect 7443 11942 7445 11994
rect 7199 11940 7205 11942
rect 7261 11940 7285 11942
rect 7341 11940 7365 11942
rect 7421 11940 7445 11942
rect 7501 11940 7507 11942
rect 7199 11931 7507 11940
rect 7576 11354 7604 12174
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7668 11014 7696 12174
rect 7748 12164 7800 12170
rect 7748 12106 7800 12112
rect 7760 11898 7788 12106
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7760 11218 7788 11834
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8036 11286 8064 11630
rect 8128 11354 8156 12242
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11898 8248 12038
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8220 11354 8248 11834
rect 8312 11642 8340 13194
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8404 12434 8432 12786
rect 8864 12782 8892 14418
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9416 14074 9444 14282
rect 9784 14074 9812 14418
rect 10060 14278 10088 14554
rect 10152 14346 10180 15030
rect 11348 14822 11376 15438
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 10265 14716 10573 14725
rect 10265 14714 10271 14716
rect 10327 14714 10351 14716
rect 10407 14714 10431 14716
rect 10487 14714 10511 14716
rect 10567 14714 10573 14716
rect 10327 14662 10329 14714
rect 10509 14662 10511 14714
rect 10265 14660 10271 14662
rect 10327 14660 10351 14662
rect 10407 14660 10431 14662
rect 10487 14660 10511 14662
rect 10567 14660 10573 14662
rect 10265 14651 10573 14660
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9048 12986 9076 13806
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8484 12640 8536 12646
rect 8536 12588 8616 12594
rect 8484 12582 8616 12588
rect 8496 12566 8616 12582
rect 8404 12406 8524 12434
rect 8496 12238 8524 12406
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8496 11898 8524 12174
rect 8588 12102 8616 12566
rect 9140 12238 9168 13806
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9232 12986 9260 13126
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9692 12238 9720 13330
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9784 12306 9812 13262
rect 10152 12918 10180 14282
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 11336 14272 11388 14278
rect 11336 14214 11388 14220
rect 10704 13938 10732 14214
rect 10925 14172 11233 14181
rect 10925 14170 10931 14172
rect 10987 14170 11011 14172
rect 11067 14170 11091 14172
rect 11147 14170 11171 14172
rect 11227 14170 11233 14172
rect 10987 14118 10989 14170
rect 11169 14118 11171 14170
rect 10925 14116 10931 14118
rect 10987 14116 11011 14118
rect 11067 14116 11091 14118
rect 11147 14116 11171 14118
rect 11227 14116 11233 14118
rect 10925 14107 11233 14116
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10265 13628 10573 13637
rect 10265 13626 10271 13628
rect 10327 13626 10351 13628
rect 10407 13626 10431 13628
rect 10487 13626 10511 13628
rect 10567 13626 10573 13628
rect 10327 13574 10329 13626
rect 10509 13574 10511 13626
rect 10265 13572 10271 13574
rect 10327 13572 10351 13574
rect 10407 13572 10431 13574
rect 10487 13572 10511 13574
rect 10567 13572 10573 13574
rect 10265 13563 10573 13572
rect 10704 13394 10732 13874
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11072 13530 11100 13806
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 11348 13462 11376 14214
rect 11440 14074 11468 15506
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11992 14958 12020 15302
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11532 14346 11560 14758
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10520 12850 10548 13262
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10612 12918 10640 13126
rect 10925 13084 11233 13093
rect 10925 13082 10931 13084
rect 10987 13082 11011 13084
rect 11067 13082 11091 13084
rect 11147 13082 11171 13084
rect 11227 13082 11233 13084
rect 10987 13030 10989 13082
rect 11169 13030 11171 13082
rect 10925 13028 10931 13030
rect 10987 13028 11011 13030
rect 11067 13028 11091 13030
rect 11147 13028 11171 13030
rect 11227 13028 11233 13030
rect 10925 13019 11233 13028
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10612 12646 10640 12854
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 9876 12442 9904 12582
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 10152 12306 10180 12582
rect 10265 12540 10573 12549
rect 10265 12538 10271 12540
rect 10327 12538 10351 12540
rect 10407 12538 10431 12540
rect 10487 12538 10511 12540
rect 10567 12538 10573 12540
rect 10327 12486 10329 12538
rect 10509 12486 10511 12538
rect 10265 12484 10271 12486
rect 10327 12484 10351 12486
rect 10407 12484 10431 12486
rect 10487 12484 10511 12486
rect 10567 12484 10573 12486
rect 10265 12475 10573 12484
rect 10704 12434 10732 12582
rect 10704 12406 10824 12434
rect 10796 12306 10824 12406
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 10152 11898 10180 12242
rect 10888 12238 10916 12582
rect 11164 12238 11192 12718
rect 11348 12714 11376 13398
rect 11440 13258 11468 14010
rect 11532 14006 11560 14282
rect 11992 14074 12020 14894
rect 12268 14618 12296 14894
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12360 14278 12388 15982
rect 12452 14414 12480 16118
rect 12912 16114 12940 16594
rect 14651 16348 14959 16357
rect 14651 16346 14657 16348
rect 14713 16346 14737 16348
rect 14793 16346 14817 16348
rect 14873 16346 14897 16348
rect 14953 16346 14959 16348
rect 14713 16294 14715 16346
rect 14895 16294 14897 16346
rect 14651 16292 14657 16294
rect 14713 16292 14737 16294
rect 14793 16292 14817 16294
rect 14873 16292 14897 16294
rect 14953 16292 14959 16294
rect 14651 16283 14959 16292
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12912 15706 12940 16050
rect 13991 15804 14299 15813
rect 13991 15802 13997 15804
rect 14053 15802 14077 15804
rect 14133 15802 14157 15804
rect 14213 15802 14237 15804
rect 14293 15802 14299 15804
rect 14053 15750 14055 15802
rect 14235 15750 14237 15802
rect 13991 15748 13997 15750
rect 14053 15748 14077 15750
rect 14133 15748 14157 15750
rect 14213 15748 14237 15750
rect 14293 15748 14299 15750
rect 13991 15739 14299 15748
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12912 15162 12940 15438
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 8312 11614 8524 11642
rect 8496 11558 8524 11614
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7199 10908 7507 10917
rect 7199 10906 7205 10908
rect 7261 10906 7285 10908
rect 7341 10906 7365 10908
rect 7421 10906 7445 10908
rect 7501 10906 7507 10908
rect 7261 10854 7263 10906
rect 7443 10854 7445 10906
rect 7199 10852 7205 10854
rect 7261 10852 7285 10854
rect 7341 10852 7365 10854
rect 7421 10852 7445 10854
rect 7501 10852 7507 10854
rect 7199 10843 7507 10852
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7208 10266 7236 10542
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7668 10130 7696 10950
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 8404 10062 8432 11086
rect 8496 11082 8524 11494
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8496 10742 8524 11018
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8588 10062 8616 11562
rect 10265 11452 10573 11461
rect 10265 11450 10271 11452
rect 10327 11450 10351 11452
rect 10407 11450 10431 11452
rect 10487 11450 10511 11452
rect 10567 11450 10573 11452
rect 10327 11398 10329 11450
rect 10509 11398 10511 11450
rect 10265 11396 10271 11398
rect 10327 11396 10351 11398
rect 10407 11396 10431 11398
rect 10487 11396 10511 11398
rect 10567 11396 10573 11398
rect 10265 11387 10573 11396
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9508 10810 9536 11086
rect 9692 10810 9720 11154
rect 10612 11014 10640 12106
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 9178 4660 9318
rect 4816 9178 4844 9454
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8634 4568 8910
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4448 8090 4476 8570
rect 4816 8362 4844 9114
rect 4908 8498 4936 9318
rect 5460 9110 5488 9522
rect 6539 9276 6847 9285
rect 6539 9274 6545 9276
rect 6601 9274 6625 9276
rect 6681 9274 6705 9276
rect 6761 9274 6785 9276
rect 6841 9274 6847 9276
rect 6601 9222 6603 9274
rect 6783 9222 6785 9274
rect 6539 9220 6545 9222
rect 6601 9220 6625 9222
rect 6681 9220 6705 9222
rect 6761 9220 6785 9222
rect 6841 9220 6847 9222
rect 6539 9211 6847 9220
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4356 7546 4384 7686
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 3896 6718 4016 6746
rect 3473 6556 3781 6565
rect 3473 6554 3479 6556
rect 3535 6554 3559 6556
rect 3615 6554 3639 6556
rect 3695 6554 3719 6556
rect 3775 6554 3781 6556
rect 3535 6502 3537 6554
rect 3717 6502 3719 6554
rect 3473 6500 3479 6502
rect 3535 6500 3559 6502
rect 3615 6500 3639 6502
rect 3695 6500 3719 6502
rect 3775 6500 3781 6502
rect 3473 6491 3781 6500
rect 3896 6458 3924 6718
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2700 5086 2820 5114
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2516 4690 2544 4966
rect 2700 4706 2728 5086
rect 2813 4924 3121 4933
rect 2813 4922 2819 4924
rect 2875 4922 2899 4924
rect 2955 4922 2979 4924
rect 3035 4922 3059 4924
rect 3115 4922 3121 4924
rect 2875 4870 2877 4922
rect 3057 4870 3059 4922
rect 2813 4868 2819 4870
rect 2875 4868 2899 4870
rect 2955 4868 2979 4870
rect 3035 4868 3059 4870
rect 3115 4868 3121 4870
rect 2813 4859 3121 4868
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 2504 4684 2556 4690
rect 2700 4678 2820 4706
rect 2504 4626 2556 4632
rect 1872 4146 1900 4626
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1872 3602 1900 4082
rect 2792 4026 2820 4678
rect 3160 4078 3188 5510
rect 3252 5030 3280 5646
rect 3344 5370 3372 5646
rect 3896 5642 3924 6394
rect 3988 6254 4016 6598
rect 4080 6322 4108 6870
rect 4172 6458 4200 6938
rect 4264 6798 4292 7142
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3988 5710 4016 6190
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3473 5468 3781 5477
rect 3473 5466 3479 5468
rect 3535 5466 3559 5468
rect 3615 5466 3639 5468
rect 3695 5466 3719 5468
rect 3775 5466 3781 5468
rect 3535 5414 3537 5466
rect 3717 5414 3719 5466
rect 3473 5412 3479 5414
rect 3535 5412 3559 5414
rect 3615 5412 3639 5414
rect 3695 5412 3719 5414
rect 3775 5412 3781 5414
rect 3473 5403 3781 5412
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3252 4146 3280 4558
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2700 3998 2820 4026
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 2700 3618 2728 3998
rect 2813 3836 3121 3845
rect 2813 3834 2819 3836
rect 2875 3834 2899 3836
rect 2955 3834 2979 3836
rect 3035 3834 3059 3836
rect 3115 3834 3121 3836
rect 2875 3782 2877 3834
rect 3057 3782 3059 3834
rect 2813 3780 2819 3782
rect 2875 3780 2899 3782
rect 2955 3780 2979 3782
rect 3035 3780 3059 3782
rect 3115 3780 3121 3782
rect 2813 3771 3121 3780
rect 1860 3596 1912 3602
rect 2700 3590 2820 3618
rect 1860 3538 1912 3544
rect 2136 3460 2188 3466
rect 2136 3402 2188 3408
rect 2148 3194 2176 3402
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2792 3058 2820 3590
rect 3252 3534 3280 4082
rect 3344 4078 3372 5102
rect 3436 4622 3464 5170
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3804 4826 3832 5102
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3473 4380 3781 4389
rect 3473 4378 3479 4380
rect 3535 4378 3559 4380
rect 3615 4378 3639 4380
rect 3695 4378 3719 4380
rect 3775 4378 3781 4380
rect 3535 4326 3537 4378
rect 3717 4326 3719 4378
rect 3473 4324 3479 4326
rect 3535 4324 3559 4326
rect 3615 4324 3639 4326
rect 3695 4324 3719 4326
rect 3775 4324 3781 4326
rect 3473 4315 3781 4324
rect 3896 4282 3924 5170
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3792 4208 3844 4214
rect 3988 4162 4016 5238
rect 4080 5166 4108 5578
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4570 4108 4966
rect 4356 4826 4384 7346
rect 5000 7342 5028 8230
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5460 7546 5488 7822
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4908 7002 4936 7210
rect 5092 7002 5120 7346
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4448 6322 4476 6666
rect 5092 6322 5120 6938
rect 5276 6934 5304 7278
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5460 6866 5488 7482
rect 6012 7206 6040 7482
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 6322 5212 6734
rect 5460 6322 5488 6802
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4344 4820 4396 4826
rect 4344 4762 4396 4768
rect 4448 4758 4476 5850
rect 4632 5370 4660 6258
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4632 4826 4660 4966
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4080 4542 4200 4570
rect 4172 4486 4200 4542
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4080 4282 4108 4422
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4172 4162 4200 4422
rect 4448 4282 4476 4694
rect 4724 4690 4752 5782
rect 5552 5778 5580 6734
rect 5644 6186 5672 6734
rect 6104 6730 6132 8366
rect 6288 7954 6316 8434
rect 6539 8188 6847 8197
rect 6539 8186 6545 8188
rect 6601 8186 6625 8188
rect 6681 8186 6705 8188
rect 6761 8186 6785 8188
rect 6841 8186 6847 8188
rect 6601 8134 6603 8186
rect 6783 8134 6785 8186
rect 6539 8132 6545 8134
rect 6601 8132 6625 8134
rect 6681 8132 6705 8134
rect 6761 8132 6785 8134
rect 6841 8132 6847 8134
rect 6539 8123 6847 8132
rect 6932 7970 6960 9930
rect 7199 9820 7507 9829
rect 7199 9818 7205 9820
rect 7261 9818 7285 9820
rect 7341 9818 7365 9820
rect 7421 9818 7445 9820
rect 7501 9818 7507 9820
rect 7261 9766 7263 9818
rect 7443 9766 7445 9818
rect 7199 9764 7205 9766
rect 7261 9764 7285 9766
rect 7341 9764 7365 9766
rect 7421 9764 7445 9766
rect 7501 9764 7507 9766
rect 7199 9755 7507 9764
rect 8220 9178 8248 9998
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8588 9110 8616 9998
rect 8758 9616 8814 9625
rect 8758 9551 8760 9560
rect 8812 9551 8814 9560
rect 8760 9522 8812 9528
rect 9232 9518 9260 10610
rect 9600 9994 9628 10610
rect 9692 10130 9720 10746
rect 10265 10364 10573 10373
rect 10265 10362 10271 10364
rect 10327 10362 10351 10364
rect 10407 10362 10431 10364
rect 10487 10362 10511 10364
rect 10567 10362 10573 10364
rect 10327 10310 10329 10362
rect 10509 10310 10511 10362
rect 10265 10308 10271 10310
rect 10327 10308 10351 10310
rect 10407 10308 10431 10310
rect 10487 10308 10511 10310
rect 10567 10308 10573 10310
rect 10265 10299 10573 10308
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9600 9704 9628 9930
rect 9600 9676 9720 9704
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 7208 8974 7236 9046
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 7196 8968 7248 8974
rect 7116 8916 7196 8922
rect 7116 8910 7248 8916
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 7116 8894 7236 8910
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6840 7942 6960 7970
rect 7024 7954 7052 8842
rect 7116 8430 7144 8894
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 7199 8732 7507 8741
rect 7199 8730 7205 8732
rect 7261 8730 7285 8732
rect 7341 8730 7365 8732
rect 7421 8730 7445 8732
rect 7501 8730 7507 8732
rect 7261 8678 7263 8730
rect 7443 8678 7445 8730
rect 7199 8676 7205 8678
rect 7261 8676 7285 8678
rect 7341 8676 7365 8678
rect 7421 8676 7445 8678
rect 7501 8676 7507 8678
rect 7199 8667 7507 8676
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7012 7948 7064 7954
rect 6288 7410 6316 7890
rect 6840 7818 6868 7942
rect 7012 7890 7064 7896
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6196 6798 6224 7142
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4908 4826 4936 5102
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 5000 4622 5028 5170
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5448 5092 5500 5098
rect 5448 5034 5500 5040
rect 5184 4826 5212 5034
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 3844 4156 4016 4162
rect 3792 4150 4016 4156
rect 3804 4134 4016 4150
rect 4080 4146 4200 4162
rect 4068 4140 4200 4146
rect 4120 4134 4200 4140
rect 4068 4082 4120 4088
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3344 3126 3372 3878
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3473 3292 3781 3301
rect 3473 3290 3479 3292
rect 3535 3290 3559 3292
rect 3615 3290 3639 3292
rect 3695 3290 3719 3292
rect 3775 3290 3781 3292
rect 3535 3238 3537 3290
rect 3717 3238 3719 3290
rect 3473 3236 3479 3238
rect 3535 3236 3559 3238
rect 3615 3236 3639 3238
rect 3695 3236 3719 3238
rect 3775 3236 3781 3238
rect 3473 3227 3781 3236
rect 3896 3194 3924 3334
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1688 2582 1716 2926
rect 4448 2854 4476 4218
rect 4632 4214 4660 4558
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4540 3738 4568 4014
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 5000 3670 5028 4558
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 5184 3398 5212 4762
rect 5460 4282 5488 5034
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4826 6040 4966
rect 6104 4826 6132 5238
rect 6196 5234 6224 5510
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6288 4690 6316 7346
rect 6539 7100 6847 7109
rect 6539 7098 6545 7100
rect 6601 7098 6625 7100
rect 6681 7098 6705 7100
rect 6761 7098 6785 7100
rect 6841 7098 6847 7100
rect 6601 7046 6603 7098
rect 6783 7046 6785 7098
rect 6539 7044 6545 7046
rect 6601 7044 6625 7046
rect 6681 7044 6705 7046
rect 6761 7044 6785 7046
rect 6841 7044 6847 7046
rect 6539 7035 6847 7044
rect 6736 6928 6788 6934
rect 6932 6916 6960 7686
rect 7116 7528 7144 8366
rect 7300 7954 7328 8570
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7300 7818 7328 7890
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7199 7644 7507 7653
rect 7199 7642 7205 7644
rect 7261 7642 7285 7644
rect 7341 7642 7365 7644
rect 7421 7642 7445 7644
rect 7501 7642 7507 7644
rect 7261 7590 7263 7642
rect 7443 7590 7445 7642
rect 7199 7588 7205 7590
rect 7261 7588 7285 7590
rect 7341 7588 7365 7590
rect 7421 7588 7445 7590
rect 7501 7588 7507 7590
rect 7199 7579 7507 7588
rect 7116 7500 7328 7528
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 6788 6888 6960 6916
rect 6736 6870 6788 6876
rect 6748 6798 6776 6870
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 7024 6730 7052 7414
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7208 7002 7236 7278
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7116 6458 7144 6802
rect 7300 6798 7328 7500
rect 7760 7478 7788 7890
rect 7944 7886 7972 8774
rect 8036 8090 8064 8910
rect 8128 8294 8156 8910
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7199 6556 7507 6565
rect 7199 6554 7205 6556
rect 7261 6554 7285 6556
rect 7341 6554 7365 6556
rect 7421 6554 7445 6556
rect 7501 6554 7507 6556
rect 7261 6502 7263 6554
rect 7443 6502 7445 6554
rect 7199 6500 7205 6502
rect 7261 6500 7285 6502
rect 7341 6500 7365 6502
rect 7421 6500 7445 6502
rect 7501 6500 7507 6502
rect 7199 6491 7507 6500
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6539 6012 6847 6021
rect 6539 6010 6545 6012
rect 6601 6010 6625 6012
rect 6681 6010 6705 6012
rect 6761 6010 6785 6012
rect 6841 6010 6847 6012
rect 6601 5958 6603 6010
rect 6783 5958 6785 6010
rect 6539 5956 6545 5958
rect 6601 5956 6625 5958
rect 6681 5956 6705 5958
rect 6761 5956 6785 5958
rect 6841 5956 6847 5958
rect 6539 5947 6847 5956
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 7012 5704 7064 5710
rect 7116 5658 7144 6054
rect 7064 5652 7144 5658
rect 7012 5646 7144 5652
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5460 3534 5488 4218
rect 5552 3738 5580 4422
rect 6104 4282 6132 4558
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6288 4146 6316 4626
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6104 3738 6132 3878
rect 6288 3738 6316 4082
rect 6472 3942 6500 5646
rect 7024 5630 7144 5646
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 5030 6868 5510
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6539 4924 6847 4933
rect 6539 4922 6545 4924
rect 6601 4922 6625 4924
rect 6681 4922 6705 4924
rect 6761 4922 6785 4924
rect 6841 4922 6847 4924
rect 6601 4870 6603 4922
rect 6783 4870 6785 4922
rect 6539 4868 6545 4870
rect 6601 4868 6625 4870
rect 6681 4868 6705 4870
rect 6761 4868 6785 4870
rect 6841 4868 6847 4870
rect 6539 4859 6847 4868
rect 7116 4808 7144 5630
rect 7199 5468 7507 5477
rect 7199 5466 7205 5468
rect 7261 5466 7285 5468
rect 7341 5466 7365 5468
rect 7421 5466 7445 5468
rect 7501 5466 7507 5468
rect 7261 5414 7263 5466
rect 7443 5414 7445 5466
rect 7199 5412 7205 5414
rect 7261 5412 7285 5414
rect 7341 5412 7365 5414
rect 7421 5412 7445 5414
rect 7501 5412 7507 5414
rect 7199 5403 7507 5412
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7576 5234 7604 5306
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7576 5030 7604 5170
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7196 4820 7248 4826
rect 7116 4780 7196 4808
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5644 3194 5672 3470
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5920 3126 5948 3470
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 6472 3058 6500 3878
rect 6539 3836 6847 3845
rect 6539 3834 6545 3836
rect 6601 3834 6625 3836
rect 6681 3834 6705 3836
rect 6761 3834 6785 3836
rect 6841 3834 6847 3836
rect 6601 3782 6603 3834
rect 6783 3782 6785 3834
rect 6539 3780 6545 3782
rect 6601 3780 6625 3782
rect 6681 3780 6705 3782
rect 6761 3780 6785 3782
rect 6841 3780 6847 3782
rect 6539 3771 6847 3780
rect 7116 3058 7144 4780
rect 7196 4762 7248 4768
rect 7199 4380 7507 4389
rect 7199 4378 7205 4380
rect 7261 4378 7285 4380
rect 7341 4378 7365 4380
rect 7421 4378 7445 4380
rect 7501 4378 7507 4380
rect 7261 4326 7263 4378
rect 7443 4326 7445 4378
rect 7199 4324 7205 4326
rect 7261 4324 7285 4326
rect 7341 4324 7365 4326
rect 7421 4324 7445 4326
rect 7501 4324 7507 4326
rect 7199 4315 7507 4324
rect 7199 3292 7507 3301
rect 7199 3290 7205 3292
rect 7261 3290 7285 3292
rect 7341 3290 7365 3292
rect 7421 3290 7445 3292
rect 7501 3290 7507 3292
rect 7261 3238 7263 3290
rect 7443 3238 7445 3290
rect 7199 3236 7205 3238
rect 7261 3236 7285 3238
rect 7341 3236 7365 3238
rect 7421 3236 7445 3238
rect 7501 3236 7507 3238
rect 7199 3227 7507 3236
rect 7576 3058 7604 4966
rect 7668 3738 7696 5034
rect 7760 4604 7788 7414
rect 7944 6866 7972 7822
rect 8128 7206 8156 8230
rect 8220 7546 8248 8978
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8312 7818 8340 8774
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8404 7546 8432 7822
rect 8208 7540 8260 7546
rect 8392 7540 8444 7546
rect 8208 7482 8260 7488
rect 8312 7500 8392 7528
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8220 7002 8248 7482
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 8312 6730 8340 7500
rect 8392 7482 8444 7488
rect 8588 7478 8616 9046
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8090 8800 8774
rect 9232 8566 9260 9454
rect 9692 9382 9720 9676
rect 10612 9674 10640 10950
rect 10796 10810 10824 12038
rect 10925 11996 11233 12005
rect 10925 11994 10931 11996
rect 10987 11994 11011 11996
rect 11067 11994 11091 11996
rect 11147 11994 11171 11996
rect 11227 11994 11233 11996
rect 10987 11942 10989 11994
rect 11169 11942 11171 11994
rect 10925 11940 10931 11942
rect 10987 11940 11011 11942
rect 11067 11940 11091 11942
rect 11147 11940 11171 11942
rect 11227 11940 11233 11942
rect 10925 11931 11233 11940
rect 11624 11626 11652 12582
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11716 12170 11744 12378
rect 11992 12306 12020 14010
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12176 12442 12204 12582
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11992 11762 12020 12242
rect 12728 12238 12756 15030
rect 13280 14822 13308 15302
rect 13268 14816 13320 14822
rect 13188 14764 13268 14770
rect 13188 14758 13320 14764
rect 13188 14742 13308 14758
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13004 14414 13032 14486
rect 13188 14414 13216 14742
rect 13464 14634 13492 15302
rect 14651 15260 14959 15269
rect 14651 15258 14657 15260
rect 14713 15258 14737 15260
rect 14793 15258 14817 15260
rect 14873 15258 14897 15260
rect 14953 15258 14959 15260
rect 14713 15206 14715 15258
rect 14895 15206 14897 15258
rect 14651 15204 14657 15206
rect 14713 15204 14737 15206
rect 14793 15204 14817 15206
rect 14873 15204 14897 15206
rect 14953 15204 14959 15206
rect 14651 15195 14959 15204
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13372 14606 13492 14634
rect 13372 14414 13400 14606
rect 13832 14482 13860 14758
rect 13991 14716 14299 14725
rect 13991 14714 13997 14716
rect 14053 14714 14077 14716
rect 14133 14714 14157 14716
rect 14213 14714 14237 14716
rect 14293 14714 14299 14716
rect 14053 14662 14055 14714
rect 14235 14662 14237 14714
rect 13991 14660 13997 14662
rect 14053 14660 14077 14662
rect 14133 14660 14157 14662
rect 14213 14660 14237 14662
rect 14293 14660 14299 14662
rect 13991 14651 14299 14660
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13004 12850 13032 14350
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13096 13530 13124 13806
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13188 12782 13216 14350
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13648 13326 13676 14214
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13924 13258 13952 14214
rect 14476 14006 14504 15098
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15304 14618 15332 14894
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14651 14172 14959 14181
rect 14651 14170 14657 14172
rect 14713 14170 14737 14172
rect 14793 14170 14817 14172
rect 14873 14170 14897 14172
rect 14953 14170 14959 14172
rect 14713 14118 14715 14170
rect 14895 14118 14897 14170
rect 14651 14116 14657 14118
rect 14713 14116 14737 14118
rect 14793 14116 14817 14118
rect 14873 14116 14897 14118
rect 14953 14116 14959 14118
rect 14651 14107 14959 14116
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 13991 13628 14299 13637
rect 13991 13626 13997 13628
rect 14053 13626 14077 13628
rect 14133 13626 14157 13628
rect 14213 13626 14237 13628
rect 14293 13626 14299 13628
rect 14053 13574 14055 13626
rect 14235 13574 14237 13626
rect 13991 13572 13997 13574
rect 14053 13572 14077 13574
rect 14133 13572 14157 13574
rect 14213 13572 14237 13574
rect 14293 13572 14299 13574
rect 13991 13563 14299 13572
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 12820 12374 12848 12718
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 12808 12368 12860 12374
rect 12808 12310 12860 12316
rect 13372 12238 13400 12582
rect 13464 12434 13492 12786
rect 13464 12406 13584 12434
rect 13556 12238 13584 12406
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 10925 10908 11233 10917
rect 10925 10906 10931 10908
rect 10987 10906 11011 10908
rect 11067 10906 11091 10908
rect 11147 10906 11171 10908
rect 11227 10906 11233 10908
rect 10987 10854 10989 10906
rect 11169 10854 11171 10906
rect 10925 10852 10931 10854
rect 10987 10852 11011 10854
rect 11067 10852 11091 10854
rect 11147 10852 11171 10854
rect 11227 10852 11233 10854
rect 10925 10843 11233 10852
rect 11348 10810 11376 11154
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11440 10674 11468 10950
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 10925 9820 11233 9829
rect 10925 9818 10931 9820
rect 10987 9818 11011 9820
rect 11067 9818 11091 9820
rect 11147 9818 11171 9820
rect 11227 9818 11233 9820
rect 10987 9766 10989 9818
rect 11169 9766 11171 9818
rect 10925 9764 10931 9766
rect 10987 9764 11011 9766
rect 11067 9764 11091 9766
rect 11147 9764 11171 9766
rect 11227 9764 11233 9766
rect 10925 9755 11233 9764
rect 11348 9722 11376 10066
rect 11532 9994 11560 11086
rect 11624 10810 11652 11562
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11716 10470 11744 11630
rect 12728 11286 12756 12174
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11898 13216 12038
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12716 11280 12768 11286
rect 12716 11222 12768 11228
rect 11796 11212 11848 11218
rect 11796 11154 11848 11160
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 11808 10674 11836 11154
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 12360 10470 12388 10950
rect 12452 10606 12480 10950
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11336 9716 11388 9722
rect 10612 9646 10824 9674
rect 11336 9658 11388 9664
rect 10796 9586 10824 9646
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10265 9276 10573 9285
rect 10265 9274 10271 9276
rect 10327 9274 10351 9276
rect 10407 9274 10431 9276
rect 10487 9274 10511 9276
rect 10567 9274 10573 9276
rect 10327 9222 10329 9274
rect 10509 9222 10511 9274
rect 10265 9220 10271 9222
rect 10327 9220 10351 9222
rect 10407 9220 10431 9222
rect 10487 9220 10511 9222
rect 10567 9220 10573 9222
rect 10265 9211 10573 9220
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9600 8634 9628 8910
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8956 7954 8984 8366
rect 9692 7954 9720 8774
rect 9784 8566 9812 8842
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8634 10272 8774
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 10265 8188 10573 8197
rect 10265 8186 10271 8188
rect 10327 8186 10351 8188
rect 10407 8186 10431 8188
rect 10487 8186 10511 8188
rect 10567 8186 10573 8188
rect 10327 8134 10329 8186
rect 10509 8134 10511 8186
rect 10265 8132 10271 8134
rect 10327 8132 10351 8134
rect 10407 8132 10431 8134
rect 10487 8132 10511 8134
rect 10567 8132 10573 8134
rect 10265 8123 10573 8132
rect 8944 7948 8996 7954
rect 8944 7890 8996 7896
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8404 6798 8432 7142
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8312 6458 8340 6666
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8588 5574 8616 6802
rect 8956 6322 8984 7890
rect 9220 7812 9272 7818
rect 9220 7754 9272 7760
rect 9232 7410 9260 7754
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 5574 8984 6258
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8312 4622 8340 5510
rect 7840 4616 7892 4622
rect 7760 4576 7840 4604
rect 7760 4146 7788 4576
rect 7840 4558 7892 4564
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8588 4486 8616 5510
rect 8956 4690 8984 5510
rect 9324 5234 9352 7142
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8312 4146 8340 4422
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7760 3534 7788 4082
rect 8588 4078 8616 4422
rect 8956 4146 8984 4626
rect 9140 4282 9168 4966
rect 9232 4690 9260 4966
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7944 3534 7972 3674
rect 8312 3534 8340 3878
rect 9508 3602 9536 4082
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 7944 3194 7972 3470
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 8312 2922 8340 3470
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 9692 2774 9720 7210
rect 10265 7100 10573 7109
rect 10265 7098 10271 7100
rect 10327 7098 10351 7100
rect 10407 7098 10431 7100
rect 10487 7098 10511 7100
rect 10567 7098 10573 7100
rect 10327 7046 10329 7098
rect 10509 7046 10511 7098
rect 10265 7044 10271 7046
rect 10327 7044 10351 7046
rect 10407 7044 10431 7046
rect 10487 7044 10511 7046
rect 10567 7044 10573 7046
rect 10265 7035 10573 7044
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9876 5914 9904 6190
rect 10265 6012 10573 6021
rect 10265 6010 10271 6012
rect 10327 6010 10351 6012
rect 10407 6010 10431 6012
rect 10487 6010 10511 6012
rect 10567 6010 10573 6012
rect 10327 5958 10329 6010
rect 10509 5958 10511 6010
rect 10265 5956 10271 5958
rect 10327 5956 10351 5958
rect 10407 5956 10431 5958
rect 10487 5956 10511 5958
rect 10567 5956 10573 5958
rect 10265 5947 10573 5956
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 10612 5710 10640 9318
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11164 8974 11192 9114
rect 11242 9072 11298 9081
rect 11242 9007 11244 9016
rect 11296 9007 11298 9016
rect 11244 8978 11296 8984
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11348 8906 11376 9522
rect 11716 9518 11744 10406
rect 12256 9716 12308 9722
rect 12256 9658 12308 9664
rect 12268 9518 12296 9658
rect 12544 9518 12572 10950
rect 12636 10538 12664 11154
rect 12820 10810 12848 11698
rect 13372 11150 13400 12174
rect 13556 11558 13584 12174
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 11286 13584 11494
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12636 10266 12664 10474
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12636 9722 12664 10202
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12820 9586 12848 10746
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11532 9110 11560 9318
rect 11520 9104 11572 9110
rect 11612 9104 11664 9110
rect 11520 9046 11572 9052
rect 11610 9072 11612 9081
rect 11664 9072 11666 9081
rect 11610 9007 11666 9016
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 10925 8732 11233 8741
rect 10925 8730 10931 8732
rect 10987 8730 11011 8732
rect 11067 8730 11091 8732
rect 11147 8730 11171 8732
rect 11227 8730 11233 8732
rect 10987 8678 10989 8730
rect 11169 8678 11171 8730
rect 10925 8676 10931 8678
rect 10987 8676 11011 8678
rect 11067 8676 11091 8678
rect 11147 8676 11171 8678
rect 11227 8676 11233 8678
rect 10925 8667 11233 8676
rect 10876 8492 10928 8498
rect 10796 8452 10876 8480
rect 10796 7750 10824 8452
rect 10876 8434 10928 8440
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 7886 11008 8230
rect 11072 8022 11100 8366
rect 11348 8294 11376 8842
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11532 8090 11560 8366
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10796 6730 10824 7686
rect 10925 7644 11233 7653
rect 10925 7642 10931 7644
rect 10987 7642 11011 7644
rect 11067 7642 11091 7644
rect 11147 7642 11171 7644
rect 11227 7642 11233 7644
rect 10987 7590 10989 7642
rect 11169 7590 11171 7642
rect 10925 7588 10931 7590
rect 10987 7588 11011 7590
rect 11067 7588 11091 7590
rect 11147 7588 11171 7590
rect 11227 7588 11233 7590
rect 10925 7579 11233 7588
rect 11348 7546 11376 7890
rect 11624 7886 11652 9007
rect 11716 8974 11744 9318
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11900 8906 11928 9318
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11716 7002 11744 7346
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 6066 10824 6666
rect 10925 6556 11233 6565
rect 10925 6554 10931 6556
rect 10987 6554 11011 6556
rect 11067 6554 11091 6556
rect 11147 6554 11171 6556
rect 11227 6554 11233 6556
rect 10987 6502 10989 6554
rect 11169 6502 11171 6554
rect 10925 6500 10931 6502
rect 10987 6500 11011 6502
rect 11067 6500 11091 6502
rect 11147 6500 11171 6502
rect 11227 6500 11233 6502
rect 10925 6491 11233 6500
rect 11532 6458 11560 6938
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10888 6066 10916 6258
rect 11716 6186 11744 6938
rect 11900 6322 11928 8842
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 10796 6038 10916 6066
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9784 3194 9812 4014
rect 9876 3738 9904 5102
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9968 3738 9996 5034
rect 10265 4924 10573 4933
rect 10265 4922 10271 4924
rect 10327 4922 10351 4924
rect 10407 4922 10431 4924
rect 10487 4922 10511 4924
rect 10567 4922 10573 4924
rect 10327 4870 10329 4922
rect 10509 4870 10511 4922
rect 10265 4868 10271 4870
rect 10327 4868 10351 4870
rect 10407 4868 10431 4870
rect 10487 4868 10511 4870
rect 10567 4868 10573 4870
rect 10265 4859 10573 4868
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 10520 4078 10548 4490
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10265 3836 10573 3845
rect 10265 3834 10271 3836
rect 10327 3834 10351 3836
rect 10407 3834 10431 3836
rect 10487 3834 10511 3836
rect 10567 3834 10573 3836
rect 10327 3782 10329 3834
rect 10509 3782 10511 3834
rect 10265 3780 10271 3782
rect 10327 3780 10351 3782
rect 10407 3780 10431 3782
rect 10487 3780 10511 3782
rect 10567 3780 10573 3782
rect 10265 3771 10573 3780
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10612 3398 10640 5170
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10704 4826 10732 5102
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10796 4706 10824 6038
rect 11992 5710 12020 8910
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8634 12204 8774
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12268 8090 12296 9046
rect 12452 8906 12480 9046
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12452 7342 12480 8842
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8498 12664 8774
rect 13464 8566 13492 11222
rect 13740 11218 13768 13126
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13832 12102 13860 12582
rect 13991 12540 14299 12549
rect 13991 12538 13997 12540
rect 14053 12538 14077 12540
rect 14133 12538 14157 12540
rect 14213 12538 14237 12540
rect 14293 12538 14299 12540
rect 14053 12486 14055 12538
rect 14235 12486 14237 12538
rect 13991 12484 13997 12486
rect 14053 12484 14077 12486
rect 14133 12484 14157 12486
rect 14213 12484 14237 12486
rect 14293 12484 14299 12486
rect 13991 12475 14299 12484
rect 14476 12434 14504 13942
rect 15028 13870 15056 14350
rect 15580 14074 15608 14894
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14568 13394 14596 13670
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12850 14596 13126
rect 14651 13084 14959 13093
rect 14651 13082 14657 13084
rect 14713 13082 14737 13084
rect 14793 13082 14817 13084
rect 14873 13082 14897 13084
rect 14953 13082 14959 13084
rect 14713 13030 14715 13082
rect 14895 13030 14897 13082
rect 14651 13028 14657 13030
rect 14713 13028 14737 13030
rect 14793 13028 14817 13030
rect 14873 13028 14897 13030
rect 14953 13028 14959 13030
rect 14651 13019 14959 13028
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14384 12406 14504 12434
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 14384 11762 14412 12406
rect 14568 12238 14596 12786
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 13991 11452 14299 11461
rect 13991 11450 13997 11452
rect 14053 11450 14077 11452
rect 14133 11450 14157 11452
rect 14213 11450 14237 11452
rect 14293 11450 14299 11452
rect 14053 11398 14055 11450
rect 14235 11398 14237 11450
rect 13991 11396 13997 11398
rect 14053 11396 14077 11398
rect 14133 11396 14157 11398
rect 14213 11396 14237 11398
rect 14293 11396 14299 11398
rect 13991 11387 14299 11396
rect 13728 11212 13780 11218
rect 13648 11172 13728 11200
rect 13648 10674 13676 11172
rect 13728 11154 13780 11160
rect 14384 11082 14412 11698
rect 14568 11694 14596 12174
rect 14651 11996 14959 12005
rect 14651 11994 14657 11996
rect 14713 11994 14737 11996
rect 14793 11994 14817 11996
rect 14873 11994 14897 11996
rect 14953 11994 14959 11996
rect 14713 11942 14715 11994
rect 14895 11942 14897 11994
rect 14651 11940 14657 11942
rect 14713 11940 14737 11942
rect 14793 11940 14817 11942
rect 14873 11940 14897 11942
rect 14953 11940 14959 11942
rect 14651 11931 14959 11940
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13648 10130 13676 10610
rect 13740 10198 13768 11018
rect 14384 10742 14412 11018
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 13991 10364 14299 10373
rect 13991 10362 13997 10364
rect 14053 10362 14077 10364
rect 14133 10362 14157 10364
rect 14213 10362 14237 10364
rect 14293 10362 14299 10364
rect 14053 10310 14055 10362
rect 14235 10310 14237 10362
rect 13991 10308 13997 10310
rect 14053 10308 14077 10310
rect 14133 10308 14157 10310
rect 14213 10308 14237 10310
rect 14293 10308 14299 10310
rect 13991 10299 14299 10308
rect 13728 10192 13780 10198
rect 13728 10134 13780 10140
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13924 9654 13952 10066
rect 14384 9654 14412 10678
rect 14476 10554 14504 10950
rect 14568 10742 14596 10950
rect 14651 10908 14959 10917
rect 14651 10906 14657 10908
rect 14713 10906 14737 10908
rect 14793 10906 14817 10908
rect 14873 10906 14897 10908
rect 14953 10906 14959 10908
rect 14713 10854 14715 10906
rect 14895 10854 14897 10906
rect 14651 10852 14657 10854
rect 14713 10852 14737 10854
rect 14793 10852 14817 10854
rect 14873 10852 14897 10854
rect 14953 10852 14959 10854
rect 14651 10843 14959 10852
rect 15028 10810 15056 11086
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14476 10526 14596 10554
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 13991 9276 14299 9285
rect 13991 9274 13997 9276
rect 14053 9274 14077 9276
rect 14133 9274 14157 9276
rect 14213 9274 14237 9276
rect 14293 9274 14299 9276
rect 14053 9222 14055 9274
rect 14235 9222 14237 9274
rect 13991 9220 13997 9222
rect 14053 9220 14077 9222
rect 14133 9220 14157 9222
rect 14213 9220 14237 9222
rect 14293 9220 14299 9222
rect 13991 9211 14299 9220
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 13464 8430 13492 8502
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 12728 7818 12756 8366
rect 13464 7886 13492 8366
rect 13832 8106 13860 8842
rect 14280 8832 14332 8838
rect 14332 8792 14412 8820
rect 14280 8774 14332 8780
rect 13991 8188 14299 8197
rect 13991 8186 13997 8188
rect 14053 8186 14077 8188
rect 14133 8186 14157 8188
rect 14213 8186 14237 8188
rect 14293 8186 14299 8188
rect 14053 8134 14055 8186
rect 14235 8134 14237 8186
rect 13991 8132 13997 8134
rect 14053 8132 14077 8134
rect 14133 8132 14157 8134
rect 14213 8132 14237 8134
rect 14293 8132 14299 8134
rect 13991 8123 14299 8132
rect 13832 8078 13952 8106
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12728 7546 12756 7754
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12728 6934 12756 7482
rect 13464 7478 13492 7822
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12084 6322 12112 6734
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6458 12204 6598
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 10925 5468 11233 5477
rect 10925 5466 10931 5468
rect 10987 5466 11011 5468
rect 11067 5466 11091 5468
rect 11147 5466 11171 5468
rect 11227 5466 11233 5468
rect 10987 5414 10989 5466
rect 11169 5414 11171 5466
rect 10925 5412 10931 5414
rect 10987 5412 11011 5414
rect 11067 5412 11091 5414
rect 11147 5412 11171 5414
rect 11227 5412 11233 5414
rect 10925 5403 11233 5412
rect 11532 5370 11560 5578
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10704 4678 10824 4706
rect 10980 4690 11008 4966
rect 10968 4684 11020 4690
rect 10704 4554 10732 4678
rect 10968 4626 11020 4632
rect 11164 4622 11192 4966
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 10612 2922 10640 3334
rect 10796 3194 10824 4558
rect 11440 4486 11468 5034
rect 11532 4758 11560 5170
rect 12084 5166 12112 6258
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12360 5710 12388 6122
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12360 5302 12388 5646
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11532 4622 11560 4694
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 10925 4380 11233 4389
rect 10925 4378 10931 4380
rect 10987 4378 11011 4380
rect 11067 4378 11091 4380
rect 11147 4378 11171 4380
rect 11227 4378 11233 4380
rect 10987 4326 10989 4378
rect 11169 4326 11171 4378
rect 10925 4324 10931 4326
rect 10987 4324 11011 4326
rect 11067 4324 11091 4326
rect 11147 4324 11171 4326
rect 11227 4324 11233 4326
rect 10925 4315 11233 4324
rect 11348 4146 11376 4422
rect 11440 4282 11468 4422
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11348 3534 11376 3946
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 10925 3292 11233 3301
rect 10925 3290 10931 3292
rect 10987 3290 11011 3292
rect 11067 3290 11091 3292
rect 11147 3290 11171 3292
rect 11227 3290 11233 3292
rect 10987 3238 10989 3290
rect 11169 3238 11171 3290
rect 10925 3236 10931 3238
rect 10987 3236 11011 3238
rect 11067 3236 11091 3238
rect 11147 3236 11171 3238
rect 11227 3236 11233 3238
rect 10925 3227 11233 3236
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 11440 3058 11468 4218
rect 11532 4078 11560 4558
rect 11612 4480 11664 4486
rect 11612 4422 11664 4428
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11532 3670 11560 4014
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11624 3058 11652 4422
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11716 3738 11744 4014
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11992 3194 12020 3470
rect 12084 3194 12112 4966
rect 12452 4486 12480 5578
rect 12636 5234 12664 5782
rect 12728 5574 12756 6870
rect 13464 6730 13492 7414
rect 13832 7002 13860 7890
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13924 6798 13952 8078
rect 14384 8022 14412 8792
rect 14476 8634 14504 8978
rect 14568 8820 14596 10526
rect 15028 10266 15056 10746
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15016 10260 15068 10266
rect 15016 10202 15068 10208
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14651 9820 14959 9829
rect 14651 9818 14657 9820
rect 14713 9818 14737 9820
rect 14793 9818 14817 9820
rect 14873 9818 14897 9820
rect 14953 9818 14959 9820
rect 14713 9766 14715 9818
rect 14895 9766 14897 9818
rect 14651 9764 14657 9766
rect 14713 9764 14737 9766
rect 14793 9764 14817 9766
rect 14873 9764 14897 9766
rect 14953 9764 14959 9766
rect 14651 9755 14959 9764
rect 15028 9178 15056 9862
rect 15120 9722 15148 10542
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15120 9058 15148 9658
rect 15396 9382 15424 11018
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 9178 15424 9318
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 14936 9042 15148 9058
rect 14924 9036 15148 9042
rect 14976 9030 15148 9036
rect 14924 8978 14976 8984
rect 14740 8832 14792 8838
rect 14568 8792 14740 8820
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8016 14424 8022
rect 14372 7958 14424 7964
rect 14476 7954 14504 8570
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14384 7478 14412 7686
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 13991 7100 14299 7109
rect 13991 7098 13997 7100
rect 14053 7098 14077 7100
rect 14133 7098 14157 7100
rect 14213 7098 14237 7100
rect 14293 7098 14299 7100
rect 14053 7046 14055 7098
rect 14235 7046 14237 7098
rect 13991 7044 13997 7046
rect 14053 7044 14077 7046
rect 14133 7044 14157 7046
rect 14213 7044 14237 7046
rect 14293 7044 14299 7046
rect 13991 7035 14299 7044
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 5370 12756 5510
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12912 5234 12940 5714
rect 13464 5370 13492 6666
rect 13991 6012 14299 6021
rect 13991 6010 13997 6012
rect 14053 6010 14077 6012
rect 14133 6010 14157 6012
rect 14213 6010 14237 6012
rect 14293 6010 14299 6012
rect 14053 5958 14055 6010
rect 14235 5958 14237 6010
rect 13991 5956 13997 5958
rect 14053 5956 14077 5958
rect 14133 5956 14157 5958
rect 14213 5956 14237 5958
rect 14293 5956 14299 5958
rect 13991 5947 14299 5956
rect 14384 5846 14412 6802
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13740 5370 13860 5386
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13728 5364 13860 5370
rect 13780 5358 13860 5364
rect 13728 5306 13780 5312
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12544 4162 12572 4966
rect 12636 4622 12664 5170
rect 12820 4826 12848 5170
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 13832 4706 13860 5358
rect 13924 4826 13952 5646
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14108 5302 14136 5510
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 13991 4924 14299 4933
rect 13991 4922 13997 4924
rect 14053 4922 14077 4924
rect 14133 4922 14157 4924
rect 14213 4922 14237 4924
rect 14293 4922 14299 4924
rect 14053 4870 14055 4922
rect 14235 4870 14237 4922
rect 13991 4868 13997 4870
rect 14053 4868 14077 4870
rect 14133 4868 14157 4870
rect 14213 4868 14237 4870
rect 14293 4868 14299 4870
rect 13991 4859 14299 4868
rect 14384 4826 14412 5782
rect 14476 5710 14504 6734
rect 14568 6662 14596 8792
rect 14740 8774 14792 8780
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14651 8732 14959 8741
rect 14651 8730 14657 8732
rect 14713 8730 14737 8732
rect 14793 8730 14817 8732
rect 14873 8730 14897 8732
rect 14953 8730 14959 8732
rect 14713 8678 14715 8730
rect 14895 8678 14897 8730
rect 14651 8676 14657 8678
rect 14713 8676 14737 8678
rect 14793 8676 14817 8678
rect 14873 8676 14897 8678
rect 14953 8676 14959 8678
rect 14651 8667 14959 8676
rect 14651 7644 14959 7653
rect 14651 7642 14657 7644
rect 14713 7642 14737 7644
rect 14793 7642 14817 7644
rect 14873 7642 14897 7644
rect 14953 7642 14959 7644
rect 14713 7590 14715 7642
rect 14895 7590 14897 7642
rect 14651 7588 14657 7590
rect 14713 7588 14737 7590
rect 14793 7588 14817 7590
rect 14873 7588 14897 7590
rect 14953 7588 14959 7590
rect 14651 7579 14959 7588
rect 15028 7410 15056 8774
rect 15396 8566 15424 9114
rect 16026 8936 16082 8945
rect 16026 8871 16028 8880
rect 16080 8871 16082 8880
rect 16028 8842 16080 8848
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15120 7546 15148 7890
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15212 7478 15240 7822
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14936 6798 14964 7278
rect 15120 7274 15148 7346
rect 15304 7342 15332 7686
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 15120 6730 15148 7210
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14651 6556 14959 6565
rect 14651 6554 14657 6556
rect 14713 6554 14737 6556
rect 14793 6554 14817 6556
rect 14873 6554 14897 6556
rect 14953 6554 14959 6556
rect 14713 6502 14715 6554
rect 14895 6502 14897 6554
rect 14651 6500 14657 6502
rect 14713 6500 14737 6502
rect 14793 6500 14817 6502
rect 14873 6500 14897 6502
rect 14953 6500 14959 6502
rect 14651 6491 14959 6500
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 14651 5468 14959 5477
rect 14651 5466 14657 5468
rect 14713 5466 14737 5468
rect 14793 5466 14817 5468
rect 14873 5466 14897 5468
rect 14953 5466 14959 5468
rect 14713 5414 14715 5466
rect 14895 5414 14897 5466
rect 14651 5412 14657 5414
rect 14713 5412 14737 5414
rect 14793 5412 14817 5414
rect 14873 5412 14897 5414
rect 14953 5412 14959 5414
rect 14651 5403 14959 5412
rect 15396 5370 15424 5646
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14292 4706 14320 4762
rect 13832 4678 13952 4706
rect 14292 4678 14596 4706
rect 12624 4616 12676 4622
rect 13832 4570 13860 4678
rect 12624 4558 12676 4564
rect 13648 4542 13860 4570
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 12728 4214 12756 4422
rect 12360 4134 12572 4162
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12624 4140 12676 4146
rect 12164 4004 12216 4010
rect 12360 3992 12388 4134
rect 12624 4082 12676 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12440 4072 12492 4078
rect 12440 4014 12492 4020
rect 12216 3964 12388 3992
rect 12164 3946 12216 3952
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 12084 2854 12112 3130
rect 12452 2854 12480 4014
rect 12636 3194 12664 4082
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 2813 2748 3121 2757
rect 2813 2746 2819 2748
rect 2875 2746 2899 2748
rect 2955 2746 2979 2748
rect 3035 2746 3059 2748
rect 3115 2746 3121 2748
rect 2875 2694 2877 2746
rect 3057 2694 3059 2746
rect 2813 2692 2819 2694
rect 2875 2692 2899 2694
rect 2955 2692 2979 2694
rect 3035 2692 3059 2694
rect 3115 2692 3121 2694
rect 2813 2683 3121 2692
rect 6539 2748 6847 2757
rect 6539 2746 6545 2748
rect 6601 2746 6625 2748
rect 6681 2746 6705 2748
rect 6761 2746 6785 2748
rect 6841 2746 6847 2748
rect 9692 2746 9904 2774
rect 6601 2694 6603 2746
rect 6783 2694 6785 2746
rect 6539 2692 6545 2694
rect 6601 2692 6625 2694
rect 6681 2692 6705 2694
rect 6761 2692 6785 2694
rect 6841 2692 6847 2694
rect 6539 2683 6847 2692
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 9876 2446 9904 2746
rect 10265 2748 10573 2757
rect 10265 2746 10271 2748
rect 10327 2746 10351 2748
rect 10407 2746 10431 2748
rect 10487 2746 10511 2748
rect 10567 2746 10573 2748
rect 10327 2694 10329 2746
rect 10509 2694 10511 2746
rect 10265 2692 10271 2694
rect 10327 2692 10351 2694
rect 10407 2692 10431 2694
rect 10487 2692 10511 2694
rect 10567 2692 10573 2694
rect 10265 2683 10573 2692
rect 12728 2446 12756 3946
rect 12820 3194 12848 4082
rect 13004 3602 13032 4082
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 13004 3058 13032 3538
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 13188 2650 13216 4422
rect 13648 3738 13676 4542
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13740 4078 13768 4422
rect 13924 4214 13952 4678
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 13728 4072 13780 4078
rect 14016 4026 14044 4558
rect 14108 4554 14320 4570
rect 14096 4548 14320 4554
rect 14148 4542 14320 4548
rect 14096 4490 14148 4496
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 4282 14228 4422
rect 14292 4282 14320 4542
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14568 4146 14596 4678
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 14651 4380 14959 4389
rect 14651 4378 14657 4380
rect 14713 4378 14737 4380
rect 14793 4378 14817 4380
rect 14873 4378 14897 4380
rect 14953 4378 14959 4380
rect 14713 4326 14715 4378
rect 14895 4326 14897 4378
rect 14651 4324 14657 4326
rect 14713 4324 14737 4326
rect 14793 4324 14817 4326
rect 14873 4324 14897 4326
rect 14953 4324 14959 4326
rect 14651 4315 14959 4324
rect 15028 4282 15056 4558
rect 15016 4276 15068 4282
rect 15016 4218 15068 4224
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 13728 4014 13780 4020
rect 13924 3998 14044 4026
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 13924 3738 13952 3998
rect 13991 3836 14299 3845
rect 13991 3834 13997 3836
rect 14053 3834 14077 3836
rect 14133 3834 14157 3836
rect 14213 3834 14237 3836
rect 14293 3834 14299 3836
rect 14053 3782 14055 3834
rect 14235 3782 14237 3834
rect 13991 3780 13997 3782
rect 14053 3780 14077 3782
rect 14133 3780 14157 3782
rect 14213 3780 14237 3782
rect 14293 3780 14299 3782
rect 13991 3771 14299 3780
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13924 2990 13952 3674
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 14016 3126 14044 3470
rect 14372 3188 14424 3194
rect 14476 3176 14504 4014
rect 14424 3148 14504 3176
rect 14372 3130 14424 3136
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 14568 2990 14596 4082
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14936 3738 14964 4014
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 15120 3534 15148 4558
rect 15476 4548 15528 4554
rect 15476 4490 15528 4496
rect 15488 4282 15516 4490
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15304 3738 15332 4014
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 14651 3292 14959 3301
rect 14651 3290 14657 3292
rect 14713 3290 14737 3292
rect 14793 3290 14817 3292
rect 14873 3290 14897 3292
rect 14953 3290 14959 3292
rect 14713 3238 14715 3290
rect 14895 3238 14897 3290
rect 14651 3236 14657 3238
rect 14713 3236 14737 3238
rect 14793 3236 14817 3238
rect 14873 3236 14897 3238
rect 14953 3236 14959 3238
rect 14651 3227 14959 3236
rect 15028 3194 15056 3402
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 13991 2748 14299 2757
rect 13991 2746 13997 2748
rect 14053 2746 14077 2748
rect 14133 2746 14157 2748
rect 14213 2746 14237 2748
rect 14293 2746 14299 2748
rect 14053 2694 14055 2746
rect 14235 2694 14237 2746
rect 13991 2692 13997 2694
rect 14053 2692 14077 2694
rect 14133 2692 14157 2694
rect 14213 2692 14237 2694
rect 14293 2692 14299 2694
rect 13991 2683 14299 2692
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 14752 2582 14780 2858
rect 15120 2854 15148 3470
rect 15672 3058 15700 4422
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 15120 2514 15148 2790
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 3473 2204 3781 2213
rect 3473 2202 3479 2204
rect 3535 2202 3559 2204
rect 3615 2202 3639 2204
rect 3695 2202 3719 2204
rect 3775 2202 3781 2204
rect 3535 2150 3537 2202
rect 3717 2150 3719 2202
rect 3473 2148 3479 2150
rect 3535 2148 3559 2150
rect 3615 2148 3639 2150
rect 3695 2148 3719 2150
rect 3775 2148 3781 2150
rect 3473 2139 3781 2148
rect 7199 2204 7507 2213
rect 7199 2202 7205 2204
rect 7261 2202 7285 2204
rect 7341 2202 7365 2204
rect 7421 2202 7445 2204
rect 7501 2202 7507 2204
rect 7261 2150 7263 2202
rect 7443 2150 7445 2202
rect 7199 2148 7205 2150
rect 7261 2148 7285 2150
rect 7341 2148 7365 2150
rect 7421 2148 7445 2150
rect 7501 2148 7507 2150
rect 7199 2139 7507 2148
rect 9692 800 9720 2246
rect 10925 2204 11233 2213
rect 10925 2202 10931 2204
rect 10987 2202 11011 2204
rect 11067 2202 11091 2204
rect 11147 2202 11171 2204
rect 11227 2202 11233 2204
rect 10987 2150 10989 2202
rect 11169 2150 11171 2202
rect 10925 2148 10931 2150
rect 10987 2148 11011 2150
rect 11067 2148 11091 2150
rect 11147 2148 11171 2150
rect 11227 2148 11233 2150
rect 10925 2139 11233 2148
rect 12912 800 12940 2246
rect 14651 2204 14959 2213
rect 14651 2202 14657 2204
rect 14713 2202 14737 2204
rect 14793 2202 14817 2204
rect 14873 2202 14897 2204
rect 14953 2202 14959 2204
rect 14713 2150 14715 2202
rect 14895 2150 14897 2202
rect 14651 2148 14657 2150
rect 14713 2148 14737 2150
rect 14793 2148 14817 2150
rect 14873 2148 14897 2150
rect 14953 2148 14959 2150
rect 14651 2139 14959 2148
rect 18 0 74 800
rect 3238 0 3294 800
rect 6458 0 6514 800
rect 9678 0 9734 800
rect 12898 0 12954 800
rect 16118 0 16174 800
<< via2 >>
rect 2819 16890 2875 16892
rect 2899 16890 2955 16892
rect 2979 16890 3035 16892
rect 3059 16890 3115 16892
rect 2819 16838 2865 16890
rect 2865 16838 2875 16890
rect 2899 16838 2929 16890
rect 2929 16838 2941 16890
rect 2941 16838 2955 16890
rect 2979 16838 2993 16890
rect 2993 16838 3005 16890
rect 3005 16838 3035 16890
rect 3059 16838 3069 16890
rect 3069 16838 3115 16890
rect 2819 16836 2875 16838
rect 2899 16836 2955 16838
rect 2979 16836 3035 16838
rect 3059 16836 3115 16838
rect 6545 16890 6601 16892
rect 6625 16890 6681 16892
rect 6705 16890 6761 16892
rect 6785 16890 6841 16892
rect 6545 16838 6591 16890
rect 6591 16838 6601 16890
rect 6625 16838 6655 16890
rect 6655 16838 6667 16890
rect 6667 16838 6681 16890
rect 6705 16838 6719 16890
rect 6719 16838 6731 16890
rect 6731 16838 6761 16890
rect 6785 16838 6795 16890
rect 6795 16838 6841 16890
rect 6545 16836 6601 16838
rect 6625 16836 6681 16838
rect 6705 16836 6761 16838
rect 6785 16836 6841 16838
rect 10271 16890 10327 16892
rect 10351 16890 10407 16892
rect 10431 16890 10487 16892
rect 10511 16890 10567 16892
rect 10271 16838 10317 16890
rect 10317 16838 10327 16890
rect 10351 16838 10381 16890
rect 10381 16838 10393 16890
rect 10393 16838 10407 16890
rect 10431 16838 10445 16890
rect 10445 16838 10457 16890
rect 10457 16838 10487 16890
rect 10511 16838 10521 16890
rect 10521 16838 10567 16890
rect 10271 16836 10327 16838
rect 10351 16836 10407 16838
rect 10431 16836 10487 16838
rect 10511 16836 10567 16838
rect 13997 16890 14053 16892
rect 14077 16890 14133 16892
rect 14157 16890 14213 16892
rect 14237 16890 14293 16892
rect 13997 16838 14043 16890
rect 14043 16838 14053 16890
rect 14077 16838 14107 16890
rect 14107 16838 14119 16890
rect 14119 16838 14133 16890
rect 14157 16838 14171 16890
rect 14171 16838 14183 16890
rect 14183 16838 14213 16890
rect 14237 16838 14247 16890
rect 14247 16838 14293 16890
rect 13997 16836 14053 16838
rect 14077 16836 14133 16838
rect 14157 16836 14213 16838
rect 14237 16836 14293 16838
rect 3479 16346 3535 16348
rect 3559 16346 3615 16348
rect 3639 16346 3695 16348
rect 3719 16346 3775 16348
rect 3479 16294 3525 16346
rect 3525 16294 3535 16346
rect 3559 16294 3589 16346
rect 3589 16294 3601 16346
rect 3601 16294 3615 16346
rect 3639 16294 3653 16346
rect 3653 16294 3665 16346
rect 3665 16294 3695 16346
rect 3719 16294 3729 16346
rect 3729 16294 3775 16346
rect 3479 16292 3535 16294
rect 3559 16292 3615 16294
rect 3639 16292 3695 16294
rect 3719 16292 3775 16294
rect 2819 15802 2875 15804
rect 2899 15802 2955 15804
rect 2979 15802 3035 15804
rect 3059 15802 3115 15804
rect 2819 15750 2865 15802
rect 2865 15750 2875 15802
rect 2899 15750 2929 15802
rect 2929 15750 2941 15802
rect 2941 15750 2955 15802
rect 2979 15750 2993 15802
rect 2993 15750 3005 15802
rect 3005 15750 3035 15802
rect 3059 15750 3069 15802
rect 3069 15750 3115 15802
rect 2819 15748 2875 15750
rect 2899 15748 2955 15750
rect 2979 15748 3035 15750
rect 3059 15748 3115 15750
rect 2819 14714 2875 14716
rect 2899 14714 2955 14716
rect 2979 14714 3035 14716
rect 3059 14714 3115 14716
rect 2819 14662 2865 14714
rect 2865 14662 2875 14714
rect 2899 14662 2929 14714
rect 2929 14662 2941 14714
rect 2941 14662 2955 14714
rect 2979 14662 2993 14714
rect 2993 14662 3005 14714
rect 3005 14662 3035 14714
rect 3059 14662 3069 14714
rect 3069 14662 3115 14714
rect 2819 14660 2875 14662
rect 2899 14660 2955 14662
rect 2979 14660 3035 14662
rect 3059 14660 3115 14662
rect 2819 13626 2875 13628
rect 2899 13626 2955 13628
rect 2979 13626 3035 13628
rect 3059 13626 3115 13628
rect 2819 13574 2865 13626
rect 2865 13574 2875 13626
rect 2899 13574 2929 13626
rect 2929 13574 2941 13626
rect 2941 13574 2955 13626
rect 2979 13574 2993 13626
rect 2993 13574 3005 13626
rect 3005 13574 3035 13626
rect 3059 13574 3069 13626
rect 3069 13574 3115 13626
rect 2819 13572 2875 13574
rect 2899 13572 2955 13574
rect 2979 13572 3035 13574
rect 3059 13572 3115 13574
rect 3479 15258 3535 15260
rect 3559 15258 3615 15260
rect 3639 15258 3695 15260
rect 3719 15258 3775 15260
rect 3479 15206 3525 15258
rect 3525 15206 3535 15258
rect 3559 15206 3589 15258
rect 3589 15206 3601 15258
rect 3601 15206 3615 15258
rect 3639 15206 3653 15258
rect 3653 15206 3665 15258
rect 3665 15206 3695 15258
rect 3719 15206 3729 15258
rect 3729 15206 3775 15258
rect 3479 15204 3535 15206
rect 3559 15204 3615 15206
rect 3639 15204 3695 15206
rect 3719 15204 3775 15206
rect 7205 16346 7261 16348
rect 7285 16346 7341 16348
rect 7365 16346 7421 16348
rect 7445 16346 7501 16348
rect 7205 16294 7251 16346
rect 7251 16294 7261 16346
rect 7285 16294 7315 16346
rect 7315 16294 7327 16346
rect 7327 16294 7341 16346
rect 7365 16294 7379 16346
rect 7379 16294 7391 16346
rect 7391 16294 7421 16346
rect 7445 16294 7455 16346
rect 7455 16294 7501 16346
rect 7205 16292 7261 16294
rect 7285 16292 7341 16294
rect 7365 16292 7421 16294
rect 7445 16292 7501 16294
rect 3479 14170 3535 14172
rect 3559 14170 3615 14172
rect 3639 14170 3695 14172
rect 3719 14170 3775 14172
rect 3479 14118 3525 14170
rect 3525 14118 3535 14170
rect 3559 14118 3589 14170
rect 3589 14118 3601 14170
rect 3601 14118 3615 14170
rect 3639 14118 3653 14170
rect 3653 14118 3665 14170
rect 3665 14118 3695 14170
rect 3719 14118 3729 14170
rect 3729 14118 3775 14170
rect 3479 14116 3535 14118
rect 3559 14116 3615 14118
rect 3639 14116 3695 14118
rect 3719 14116 3775 14118
rect 2819 12538 2875 12540
rect 2899 12538 2955 12540
rect 2979 12538 3035 12540
rect 3059 12538 3115 12540
rect 2819 12486 2865 12538
rect 2865 12486 2875 12538
rect 2899 12486 2929 12538
rect 2929 12486 2941 12538
rect 2941 12486 2955 12538
rect 2979 12486 2993 12538
rect 2993 12486 3005 12538
rect 3005 12486 3035 12538
rect 3059 12486 3069 12538
rect 3069 12486 3115 12538
rect 2819 12484 2875 12486
rect 2899 12484 2955 12486
rect 2979 12484 3035 12486
rect 3059 12484 3115 12486
rect 3479 13082 3535 13084
rect 3559 13082 3615 13084
rect 3639 13082 3695 13084
rect 3719 13082 3775 13084
rect 3479 13030 3525 13082
rect 3525 13030 3535 13082
rect 3559 13030 3589 13082
rect 3589 13030 3601 13082
rect 3601 13030 3615 13082
rect 3639 13030 3653 13082
rect 3653 13030 3665 13082
rect 3665 13030 3695 13082
rect 3719 13030 3729 13082
rect 3729 13030 3775 13082
rect 3479 13028 3535 13030
rect 3559 13028 3615 13030
rect 3639 13028 3695 13030
rect 3719 13028 3775 13030
rect 3479 11994 3535 11996
rect 3559 11994 3615 11996
rect 3639 11994 3695 11996
rect 3719 11994 3775 11996
rect 3479 11942 3525 11994
rect 3525 11942 3535 11994
rect 3559 11942 3589 11994
rect 3589 11942 3601 11994
rect 3601 11942 3615 11994
rect 3639 11942 3653 11994
rect 3653 11942 3665 11994
rect 3665 11942 3695 11994
rect 3719 11942 3729 11994
rect 3729 11942 3775 11994
rect 3479 11940 3535 11942
rect 3559 11940 3615 11942
rect 3639 11940 3695 11942
rect 3719 11940 3775 11942
rect 2819 11450 2875 11452
rect 2899 11450 2955 11452
rect 2979 11450 3035 11452
rect 3059 11450 3115 11452
rect 2819 11398 2865 11450
rect 2865 11398 2875 11450
rect 2899 11398 2929 11450
rect 2929 11398 2941 11450
rect 2941 11398 2955 11450
rect 2979 11398 2993 11450
rect 2993 11398 3005 11450
rect 3005 11398 3035 11450
rect 3059 11398 3069 11450
rect 3069 11398 3115 11450
rect 2819 11396 2875 11398
rect 2899 11396 2955 11398
rect 2979 11396 3035 11398
rect 3059 11396 3115 11398
rect 938 10240 994 10296
rect 2819 10362 2875 10364
rect 2899 10362 2955 10364
rect 2979 10362 3035 10364
rect 3059 10362 3115 10364
rect 2819 10310 2865 10362
rect 2865 10310 2875 10362
rect 2899 10310 2929 10362
rect 2929 10310 2941 10362
rect 2941 10310 2955 10362
rect 2979 10310 2993 10362
rect 2993 10310 3005 10362
rect 3005 10310 3035 10362
rect 3059 10310 3069 10362
rect 3069 10310 3115 10362
rect 2819 10308 2875 10310
rect 2899 10308 2955 10310
rect 2979 10308 3035 10310
rect 3059 10308 3115 10310
rect 6545 15802 6601 15804
rect 6625 15802 6681 15804
rect 6705 15802 6761 15804
rect 6785 15802 6841 15804
rect 6545 15750 6591 15802
rect 6591 15750 6601 15802
rect 6625 15750 6655 15802
rect 6655 15750 6667 15802
rect 6667 15750 6681 15802
rect 6705 15750 6719 15802
rect 6719 15750 6731 15802
rect 6731 15750 6761 15802
rect 6785 15750 6795 15802
rect 6795 15750 6841 15802
rect 6545 15748 6601 15750
rect 6625 15748 6681 15750
rect 6705 15748 6761 15750
rect 6785 15748 6841 15750
rect 6545 14714 6601 14716
rect 6625 14714 6681 14716
rect 6705 14714 6761 14716
rect 6785 14714 6841 14716
rect 6545 14662 6591 14714
rect 6591 14662 6601 14714
rect 6625 14662 6655 14714
rect 6655 14662 6667 14714
rect 6667 14662 6681 14714
rect 6705 14662 6719 14714
rect 6719 14662 6731 14714
rect 6731 14662 6761 14714
rect 6785 14662 6795 14714
rect 6795 14662 6841 14714
rect 6545 14660 6601 14662
rect 6625 14660 6681 14662
rect 6705 14660 6761 14662
rect 6785 14660 6841 14662
rect 6545 13626 6601 13628
rect 6625 13626 6681 13628
rect 6705 13626 6761 13628
rect 6785 13626 6841 13628
rect 6545 13574 6591 13626
rect 6591 13574 6601 13626
rect 6625 13574 6655 13626
rect 6655 13574 6667 13626
rect 6667 13574 6681 13626
rect 6705 13574 6719 13626
rect 6719 13574 6731 13626
rect 6731 13574 6761 13626
rect 6785 13574 6795 13626
rect 6795 13574 6841 13626
rect 6545 13572 6601 13574
rect 6625 13572 6681 13574
rect 6705 13572 6761 13574
rect 6785 13572 6841 13574
rect 7205 15258 7261 15260
rect 7285 15258 7341 15260
rect 7365 15258 7421 15260
rect 7445 15258 7501 15260
rect 7205 15206 7251 15258
rect 7251 15206 7261 15258
rect 7285 15206 7315 15258
rect 7315 15206 7327 15258
rect 7327 15206 7341 15258
rect 7365 15206 7379 15258
rect 7379 15206 7391 15258
rect 7391 15206 7421 15258
rect 7445 15206 7455 15258
rect 7455 15206 7501 15258
rect 7205 15204 7261 15206
rect 7285 15204 7341 15206
rect 7365 15204 7421 15206
rect 7445 15204 7501 15206
rect 10931 16346 10987 16348
rect 11011 16346 11067 16348
rect 11091 16346 11147 16348
rect 11171 16346 11227 16348
rect 10931 16294 10977 16346
rect 10977 16294 10987 16346
rect 11011 16294 11041 16346
rect 11041 16294 11053 16346
rect 11053 16294 11067 16346
rect 11091 16294 11105 16346
rect 11105 16294 11117 16346
rect 11117 16294 11147 16346
rect 11171 16294 11181 16346
rect 11181 16294 11227 16346
rect 10931 16292 10987 16294
rect 11011 16292 11067 16294
rect 11091 16292 11147 16294
rect 11171 16292 11227 16294
rect 10271 15802 10327 15804
rect 10351 15802 10407 15804
rect 10431 15802 10487 15804
rect 10511 15802 10567 15804
rect 10271 15750 10317 15802
rect 10317 15750 10327 15802
rect 10351 15750 10381 15802
rect 10381 15750 10393 15802
rect 10393 15750 10407 15802
rect 10431 15750 10445 15802
rect 10445 15750 10457 15802
rect 10457 15750 10487 15802
rect 10511 15750 10521 15802
rect 10521 15750 10567 15802
rect 10271 15748 10327 15750
rect 10351 15748 10407 15750
rect 10431 15748 10487 15750
rect 10511 15748 10567 15750
rect 10931 15258 10987 15260
rect 11011 15258 11067 15260
rect 11091 15258 11147 15260
rect 11171 15258 11227 15260
rect 10931 15206 10977 15258
rect 10977 15206 10987 15258
rect 11011 15206 11041 15258
rect 11041 15206 11053 15258
rect 11053 15206 11067 15258
rect 11091 15206 11105 15258
rect 11105 15206 11117 15258
rect 11117 15206 11147 15258
rect 11171 15206 11181 15258
rect 11181 15206 11227 15258
rect 10931 15204 10987 15206
rect 11011 15204 11067 15206
rect 11091 15204 11147 15206
rect 11171 15204 11227 15206
rect 6545 12538 6601 12540
rect 6625 12538 6681 12540
rect 6705 12538 6761 12540
rect 6785 12538 6841 12540
rect 6545 12486 6591 12538
rect 6591 12486 6601 12538
rect 6625 12486 6655 12538
rect 6655 12486 6667 12538
rect 6667 12486 6681 12538
rect 6705 12486 6719 12538
rect 6719 12486 6731 12538
rect 6731 12486 6761 12538
rect 6785 12486 6795 12538
rect 6795 12486 6841 12538
rect 6545 12484 6601 12486
rect 6625 12484 6681 12486
rect 6705 12484 6761 12486
rect 6785 12484 6841 12486
rect 7205 14170 7261 14172
rect 7285 14170 7341 14172
rect 7365 14170 7421 14172
rect 7445 14170 7501 14172
rect 7205 14118 7251 14170
rect 7251 14118 7261 14170
rect 7285 14118 7315 14170
rect 7315 14118 7327 14170
rect 7327 14118 7341 14170
rect 7365 14118 7379 14170
rect 7379 14118 7391 14170
rect 7391 14118 7421 14170
rect 7445 14118 7455 14170
rect 7455 14118 7501 14170
rect 7205 14116 7261 14118
rect 7285 14116 7341 14118
rect 7365 14116 7421 14118
rect 7445 14116 7501 14118
rect 7205 13082 7261 13084
rect 7285 13082 7341 13084
rect 7365 13082 7421 13084
rect 7445 13082 7501 13084
rect 7205 13030 7251 13082
rect 7251 13030 7261 13082
rect 7285 13030 7315 13082
rect 7315 13030 7327 13082
rect 7327 13030 7341 13082
rect 7365 13030 7379 13082
rect 7379 13030 7391 13082
rect 7391 13030 7421 13082
rect 7445 13030 7455 13082
rect 7455 13030 7501 13082
rect 7205 13028 7261 13030
rect 7285 13028 7341 13030
rect 7365 13028 7421 13030
rect 7445 13028 7501 13030
rect 6545 11450 6601 11452
rect 6625 11450 6681 11452
rect 6705 11450 6761 11452
rect 6785 11450 6841 11452
rect 6545 11398 6591 11450
rect 6591 11398 6601 11450
rect 6625 11398 6655 11450
rect 6655 11398 6667 11450
rect 6667 11398 6681 11450
rect 6705 11398 6719 11450
rect 6719 11398 6731 11450
rect 6731 11398 6761 11450
rect 6785 11398 6795 11450
rect 6795 11398 6841 11450
rect 6545 11396 6601 11398
rect 6625 11396 6681 11398
rect 6705 11396 6761 11398
rect 6785 11396 6841 11398
rect 3479 10906 3535 10908
rect 3559 10906 3615 10908
rect 3639 10906 3695 10908
rect 3719 10906 3775 10908
rect 3479 10854 3525 10906
rect 3525 10854 3535 10906
rect 3559 10854 3589 10906
rect 3589 10854 3601 10906
rect 3601 10854 3615 10906
rect 3639 10854 3653 10906
rect 3653 10854 3665 10906
rect 3665 10854 3695 10906
rect 3719 10854 3729 10906
rect 3729 10854 3775 10906
rect 3479 10852 3535 10854
rect 3559 10852 3615 10854
rect 3639 10852 3695 10854
rect 3719 10852 3775 10854
rect 3479 9818 3535 9820
rect 3559 9818 3615 9820
rect 3639 9818 3695 9820
rect 3719 9818 3775 9820
rect 3479 9766 3525 9818
rect 3525 9766 3535 9818
rect 3559 9766 3589 9818
rect 3589 9766 3601 9818
rect 3601 9766 3615 9818
rect 3639 9766 3653 9818
rect 3653 9766 3665 9818
rect 3665 9766 3695 9818
rect 3719 9766 3729 9818
rect 3729 9766 3775 9818
rect 3479 9764 3535 9766
rect 3559 9764 3615 9766
rect 3639 9764 3695 9766
rect 3719 9764 3775 9766
rect 662 9560 718 9616
rect 2819 9274 2875 9276
rect 2899 9274 2955 9276
rect 2979 9274 3035 9276
rect 3059 9274 3115 9276
rect 2819 9222 2865 9274
rect 2865 9222 2875 9274
rect 2899 9222 2929 9274
rect 2929 9222 2941 9274
rect 2941 9222 2955 9274
rect 2979 9222 2993 9274
rect 2993 9222 3005 9274
rect 3005 9222 3035 9274
rect 3059 9222 3069 9274
rect 3069 9222 3115 9274
rect 2819 9220 2875 9222
rect 2899 9220 2955 9222
rect 2979 9220 3035 9222
rect 3059 9220 3115 9222
rect 2819 8186 2875 8188
rect 2899 8186 2955 8188
rect 2979 8186 3035 8188
rect 3059 8186 3115 8188
rect 2819 8134 2865 8186
rect 2865 8134 2875 8186
rect 2899 8134 2929 8186
rect 2929 8134 2941 8186
rect 2941 8134 2955 8186
rect 2979 8134 2993 8186
rect 2993 8134 3005 8186
rect 3005 8134 3035 8186
rect 3059 8134 3069 8186
rect 3069 8134 3115 8186
rect 2819 8132 2875 8134
rect 2899 8132 2955 8134
rect 2979 8132 3035 8134
rect 3059 8132 3115 8134
rect 2819 7098 2875 7100
rect 2899 7098 2955 7100
rect 2979 7098 3035 7100
rect 3059 7098 3115 7100
rect 2819 7046 2865 7098
rect 2865 7046 2875 7098
rect 2899 7046 2929 7098
rect 2929 7046 2941 7098
rect 2941 7046 2955 7098
rect 2979 7046 2993 7098
rect 2993 7046 3005 7098
rect 3005 7046 3035 7098
rect 3059 7046 3069 7098
rect 3069 7046 3115 7098
rect 2819 7044 2875 7046
rect 2899 7044 2955 7046
rect 2979 7044 3035 7046
rect 3059 7044 3115 7046
rect 3479 8730 3535 8732
rect 3559 8730 3615 8732
rect 3639 8730 3695 8732
rect 3719 8730 3775 8732
rect 3479 8678 3525 8730
rect 3525 8678 3535 8730
rect 3559 8678 3589 8730
rect 3589 8678 3601 8730
rect 3601 8678 3615 8730
rect 3639 8678 3653 8730
rect 3653 8678 3665 8730
rect 3665 8678 3695 8730
rect 3719 8678 3729 8730
rect 3729 8678 3775 8730
rect 3479 8676 3535 8678
rect 3559 8676 3615 8678
rect 3639 8676 3695 8678
rect 3719 8676 3775 8678
rect 3479 7642 3535 7644
rect 3559 7642 3615 7644
rect 3639 7642 3695 7644
rect 3719 7642 3775 7644
rect 3479 7590 3525 7642
rect 3525 7590 3535 7642
rect 3559 7590 3589 7642
rect 3589 7590 3601 7642
rect 3601 7590 3615 7642
rect 3639 7590 3653 7642
rect 3653 7590 3665 7642
rect 3665 7590 3695 7642
rect 3719 7590 3729 7642
rect 3729 7590 3775 7642
rect 3479 7588 3535 7590
rect 3559 7588 3615 7590
rect 3639 7588 3695 7590
rect 3719 7588 3775 7590
rect 2819 6010 2875 6012
rect 2899 6010 2955 6012
rect 2979 6010 3035 6012
rect 3059 6010 3115 6012
rect 2819 5958 2865 6010
rect 2865 5958 2875 6010
rect 2899 5958 2929 6010
rect 2929 5958 2941 6010
rect 2941 5958 2955 6010
rect 2979 5958 2993 6010
rect 2993 5958 3005 6010
rect 3005 5958 3035 6010
rect 3059 5958 3069 6010
rect 3069 5958 3115 6010
rect 2819 5956 2875 5958
rect 2899 5956 2955 5958
rect 2979 5956 3035 5958
rect 3059 5956 3115 5958
rect 6545 10362 6601 10364
rect 6625 10362 6681 10364
rect 6705 10362 6761 10364
rect 6785 10362 6841 10364
rect 6545 10310 6591 10362
rect 6591 10310 6601 10362
rect 6625 10310 6655 10362
rect 6655 10310 6667 10362
rect 6667 10310 6681 10362
rect 6705 10310 6719 10362
rect 6719 10310 6731 10362
rect 6731 10310 6761 10362
rect 6785 10310 6795 10362
rect 6795 10310 6841 10362
rect 6545 10308 6601 10310
rect 6625 10308 6681 10310
rect 6705 10308 6761 10310
rect 6785 10308 6841 10310
rect 7205 11994 7261 11996
rect 7285 11994 7341 11996
rect 7365 11994 7421 11996
rect 7445 11994 7501 11996
rect 7205 11942 7251 11994
rect 7251 11942 7261 11994
rect 7285 11942 7315 11994
rect 7315 11942 7327 11994
rect 7327 11942 7341 11994
rect 7365 11942 7379 11994
rect 7379 11942 7391 11994
rect 7391 11942 7421 11994
rect 7445 11942 7455 11994
rect 7455 11942 7501 11994
rect 7205 11940 7261 11942
rect 7285 11940 7341 11942
rect 7365 11940 7421 11942
rect 7445 11940 7501 11942
rect 10271 14714 10327 14716
rect 10351 14714 10407 14716
rect 10431 14714 10487 14716
rect 10511 14714 10567 14716
rect 10271 14662 10317 14714
rect 10317 14662 10327 14714
rect 10351 14662 10381 14714
rect 10381 14662 10393 14714
rect 10393 14662 10407 14714
rect 10431 14662 10445 14714
rect 10445 14662 10457 14714
rect 10457 14662 10487 14714
rect 10511 14662 10521 14714
rect 10521 14662 10567 14714
rect 10271 14660 10327 14662
rect 10351 14660 10407 14662
rect 10431 14660 10487 14662
rect 10511 14660 10567 14662
rect 10931 14170 10987 14172
rect 11011 14170 11067 14172
rect 11091 14170 11147 14172
rect 11171 14170 11227 14172
rect 10931 14118 10977 14170
rect 10977 14118 10987 14170
rect 11011 14118 11041 14170
rect 11041 14118 11053 14170
rect 11053 14118 11067 14170
rect 11091 14118 11105 14170
rect 11105 14118 11117 14170
rect 11117 14118 11147 14170
rect 11171 14118 11181 14170
rect 11181 14118 11227 14170
rect 10931 14116 10987 14118
rect 11011 14116 11067 14118
rect 11091 14116 11147 14118
rect 11171 14116 11227 14118
rect 10271 13626 10327 13628
rect 10351 13626 10407 13628
rect 10431 13626 10487 13628
rect 10511 13626 10567 13628
rect 10271 13574 10317 13626
rect 10317 13574 10327 13626
rect 10351 13574 10381 13626
rect 10381 13574 10393 13626
rect 10393 13574 10407 13626
rect 10431 13574 10445 13626
rect 10445 13574 10457 13626
rect 10457 13574 10487 13626
rect 10511 13574 10521 13626
rect 10521 13574 10567 13626
rect 10271 13572 10327 13574
rect 10351 13572 10407 13574
rect 10431 13572 10487 13574
rect 10511 13572 10567 13574
rect 10931 13082 10987 13084
rect 11011 13082 11067 13084
rect 11091 13082 11147 13084
rect 11171 13082 11227 13084
rect 10931 13030 10977 13082
rect 10977 13030 10987 13082
rect 11011 13030 11041 13082
rect 11041 13030 11053 13082
rect 11053 13030 11067 13082
rect 11091 13030 11105 13082
rect 11105 13030 11117 13082
rect 11117 13030 11147 13082
rect 11171 13030 11181 13082
rect 11181 13030 11227 13082
rect 10931 13028 10987 13030
rect 11011 13028 11067 13030
rect 11091 13028 11147 13030
rect 11171 13028 11227 13030
rect 10271 12538 10327 12540
rect 10351 12538 10407 12540
rect 10431 12538 10487 12540
rect 10511 12538 10567 12540
rect 10271 12486 10317 12538
rect 10317 12486 10327 12538
rect 10351 12486 10381 12538
rect 10381 12486 10393 12538
rect 10393 12486 10407 12538
rect 10431 12486 10445 12538
rect 10445 12486 10457 12538
rect 10457 12486 10487 12538
rect 10511 12486 10521 12538
rect 10521 12486 10567 12538
rect 10271 12484 10327 12486
rect 10351 12484 10407 12486
rect 10431 12484 10487 12486
rect 10511 12484 10567 12486
rect 14657 16346 14713 16348
rect 14737 16346 14793 16348
rect 14817 16346 14873 16348
rect 14897 16346 14953 16348
rect 14657 16294 14703 16346
rect 14703 16294 14713 16346
rect 14737 16294 14767 16346
rect 14767 16294 14779 16346
rect 14779 16294 14793 16346
rect 14817 16294 14831 16346
rect 14831 16294 14843 16346
rect 14843 16294 14873 16346
rect 14897 16294 14907 16346
rect 14907 16294 14953 16346
rect 14657 16292 14713 16294
rect 14737 16292 14793 16294
rect 14817 16292 14873 16294
rect 14897 16292 14953 16294
rect 13997 15802 14053 15804
rect 14077 15802 14133 15804
rect 14157 15802 14213 15804
rect 14237 15802 14293 15804
rect 13997 15750 14043 15802
rect 14043 15750 14053 15802
rect 14077 15750 14107 15802
rect 14107 15750 14119 15802
rect 14119 15750 14133 15802
rect 14157 15750 14171 15802
rect 14171 15750 14183 15802
rect 14183 15750 14213 15802
rect 14237 15750 14247 15802
rect 14247 15750 14293 15802
rect 13997 15748 14053 15750
rect 14077 15748 14133 15750
rect 14157 15748 14213 15750
rect 14237 15748 14293 15750
rect 7205 10906 7261 10908
rect 7285 10906 7341 10908
rect 7365 10906 7421 10908
rect 7445 10906 7501 10908
rect 7205 10854 7251 10906
rect 7251 10854 7261 10906
rect 7285 10854 7315 10906
rect 7315 10854 7327 10906
rect 7327 10854 7341 10906
rect 7365 10854 7379 10906
rect 7379 10854 7391 10906
rect 7391 10854 7421 10906
rect 7445 10854 7455 10906
rect 7455 10854 7501 10906
rect 7205 10852 7261 10854
rect 7285 10852 7341 10854
rect 7365 10852 7421 10854
rect 7445 10852 7501 10854
rect 10271 11450 10327 11452
rect 10351 11450 10407 11452
rect 10431 11450 10487 11452
rect 10511 11450 10567 11452
rect 10271 11398 10317 11450
rect 10317 11398 10327 11450
rect 10351 11398 10381 11450
rect 10381 11398 10393 11450
rect 10393 11398 10407 11450
rect 10431 11398 10445 11450
rect 10445 11398 10457 11450
rect 10457 11398 10487 11450
rect 10511 11398 10521 11450
rect 10521 11398 10567 11450
rect 10271 11396 10327 11398
rect 10351 11396 10407 11398
rect 10431 11396 10487 11398
rect 10511 11396 10567 11398
rect 6545 9274 6601 9276
rect 6625 9274 6681 9276
rect 6705 9274 6761 9276
rect 6785 9274 6841 9276
rect 6545 9222 6591 9274
rect 6591 9222 6601 9274
rect 6625 9222 6655 9274
rect 6655 9222 6667 9274
rect 6667 9222 6681 9274
rect 6705 9222 6719 9274
rect 6719 9222 6731 9274
rect 6731 9222 6761 9274
rect 6785 9222 6795 9274
rect 6795 9222 6841 9274
rect 6545 9220 6601 9222
rect 6625 9220 6681 9222
rect 6705 9220 6761 9222
rect 6785 9220 6841 9222
rect 3479 6554 3535 6556
rect 3559 6554 3615 6556
rect 3639 6554 3695 6556
rect 3719 6554 3775 6556
rect 3479 6502 3525 6554
rect 3525 6502 3535 6554
rect 3559 6502 3589 6554
rect 3589 6502 3601 6554
rect 3601 6502 3615 6554
rect 3639 6502 3653 6554
rect 3653 6502 3665 6554
rect 3665 6502 3695 6554
rect 3719 6502 3729 6554
rect 3729 6502 3775 6554
rect 3479 6500 3535 6502
rect 3559 6500 3615 6502
rect 3639 6500 3695 6502
rect 3719 6500 3775 6502
rect 2819 4922 2875 4924
rect 2899 4922 2955 4924
rect 2979 4922 3035 4924
rect 3059 4922 3115 4924
rect 2819 4870 2865 4922
rect 2865 4870 2875 4922
rect 2899 4870 2929 4922
rect 2929 4870 2941 4922
rect 2941 4870 2955 4922
rect 2979 4870 2993 4922
rect 2993 4870 3005 4922
rect 3005 4870 3035 4922
rect 3059 4870 3069 4922
rect 3069 4870 3115 4922
rect 2819 4868 2875 4870
rect 2899 4868 2955 4870
rect 2979 4868 3035 4870
rect 3059 4868 3115 4870
rect 3479 5466 3535 5468
rect 3559 5466 3615 5468
rect 3639 5466 3695 5468
rect 3719 5466 3775 5468
rect 3479 5414 3525 5466
rect 3525 5414 3535 5466
rect 3559 5414 3589 5466
rect 3589 5414 3601 5466
rect 3601 5414 3615 5466
rect 3639 5414 3653 5466
rect 3653 5414 3665 5466
rect 3665 5414 3695 5466
rect 3719 5414 3729 5466
rect 3729 5414 3775 5466
rect 3479 5412 3535 5414
rect 3559 5412 3615 5414
rect 3639 5412 3695 5414
rect 3719 5412 3775 5414
rect 2819 3834 2875 3836
rect 2899 3834 2955 3836
rect 2979 3834 3035 3836
rect 3059 3834 3115 3836
rect 2819 3782 2865 3834
rect 2865 3782 2875 3834
rect 2899 3782 2929 3834
rect 2929 3782 2941 3834
rect 2941 3782 2955 3834
rect 2979 3782 2993 3834
rect 2993 3782 3005 3834
rect 3005 3782 3035 3834
rect 3059 3782 3069 3834
rect 3069 3782 3115 3834
rect 2819 3780 2875 3782
rect 2899 3780 2955 3782
rect 2979 3780 3035 3782
rect 3059 3780 3115 3782
rect 3479 4378 3535 4380
rect 3559 4378 3615 4380
rect 3639 4378 3695 4380
rect 3719 4378 3775 4380
rect 3479 4326 3525 4378
rect 3525 4326 3535 4378
rect 3559 4326 3589 4378
rect 3589 4326 3601 4378
rect 3601 4326 3615 4378
rect 3639 4326 3653 4378
rect 3653 4326 3665 4378
rect 3665 4326 3695 4378
rect 3719 4326 3729 4378
rect 3729 4326 3775 4378
rect 3479 4324 3535 4326
rect 3559 4324 3615 4326
rect 3639 4324 3695 4326
rect 3719 4324 3775 4326
rect 6545 8186 6601 8188
rect 6625 8186 6681 8188
rect 6705 8186 6761 8188
rect 6785 8186 6841 8188
rect 6545 8134 6591 8186
rect 6591 8134 6601 8186
rect 6625 8134 6655 8186
rect 6655 8134 6667 8186
rect 6667 8134 6681 8186
rect 6705 8134 6719 8186
rect 6719 8134 6731 8186
rect 6731 8134 6761 8186
rect 6785 8134 6795 8186
rect 6795 8134 6841 8186
rect 6545 8132 6601 8134
rect 6625 8132 6681 8134
rect 6705 8132 6761 8134
rect 6785 8132 6841 8134
rect 7205 9818 7261 9820
rect 7285 9818 7341 9820
rect 7365 9818 7421 9820
rect 7445 9818 7501 9820
rect 7205 9766 7251 9818
rect 7251 9766 7261 9818
rect 7285 9766 7315 9818
rect 7315 9766 7327 9818
rect 7327 9766 7341 9818
rect 7365 9766 7379 9818
rect 7379 9766 7391 9818
rect 7391 9766 7421 9818
rect 7445 9766 7455 9818
rect 7455 9766 7501 9818
rect 7205 9764 7261 9766
rect 7285 9764 7341 9766
rect 7365 9764 7421 9766
rect 7445 9764 7501 9766
rect 8758 9580 8814 9616
rect 8758 9560 8760 9580
rect 8760 9560 8812 9580
rect 8812 9560 8814 9580
rect 10271 10362 10327 10364
rect 10351 10362 10407 10364
rect 10431 10362 10487 10364
rect 10511 10362 10567 10364
rect 10271 10310 10317 10362
rect 10317 10310 10327 10362
rect 10351 10310 10381 10362
rect 10381 10310 10393 10362
rect 10393 10310 10407 10362
rect 10431 10310 10445 10362
rect 10445 10310 10457 10362
rect 10457 10310 10487 10362
rect 10511 10310 10521 10362
rect 10521 10310 10567 10362
rect 10271 10308 10327 10310
rect 10351 10308 10407 10310
rect 10431 10308 10487 10310
rect 10511 10308 10567 10310
rect 7205 8730 7261 8732
rect 7285 8730 7341 8732
rect 7365 8730 7421 8732
rect 7445 8730 7501 8732
rect 7205 8678 7251 8730
rect 7251 8678 7261 8730
rect 7285 8678 7315 8730
rect 7315 8678 7327 8730
rect 7327 8678 7341 8730
rect 7365 8678 7379 8730
rect 7379 8678 7391 8730
rect 7391 8678 7421 8730
rect 7445 8678 7455 8730
rect 7455 8678 7501 8730
rect 7205 8676 7261 8678
rect 7285 8676 7341 8678
rect 7365 8676 7421 8678
rect 7445 8676 7501 8678
rect 3479 3290 3535 3292
rect 3559 3290 3615 3292
rect 3639 3290 3695 3292
rect 3719 3290 3775 3292
rect 3479 3238 3525 3290
rect 3525 3238 3535 3290
rect 3559 3238 3589 3290
rect 3589 3238 3601 3290
rect 3601 3238 3615 3290
rect 3639 3238 3653 3290
rect 3653 3238 3665 3290
rect 3665 3238 3695 3290
rect 3719 3238 3729 3290
rect 3729 3238 3775 3290
rect 3479 3236 3535 3238
rect 3559 3236 3615 3238
rect 3639 3236 3695 3238
rect 3719 3236 3775 3238
rect 6545 7098 6601 7100
rect 6625 7098 6681 7100
rect 6705 7098 6761 7100
rect 6785 7098 6841 7100
rect 6545 7046 6591 7098
rect 6591 7046 6601 7098
rect 6625 7046 6655 7098
rect 6655 7046 6667 7098
rect 6667 7046 6681 7098
rect 6705 7046 6719 7098
rect 6719 7046 6731 7098
rect 6731 7046 6761 7098
rect 6785 7046 6795 7098
rect 6795 7046 6841 7098
rect 6545 7044 6601 7046
rect 6625 7044 6681 7046
rect 6705 7044 6761 7046
rect 6785 7044 6841 7046
rect 7205 7642 7261 7644
rect 7285 7642 7341 7644
rect 7365 7642 7421 7644
rect 7445 7642 7501 7644
rect 7205 7590 7251 7642
rect 7251 7590 7261 7642
rect 7285 7590 7315 7642
rect 7315 7590 7327 7642
rect 7327 7590 7341 7642
rect 7365 7590 7379 7642
rect 7379 7590 7391 7642
rect 7391 7590 7421 7642
rect 7445 7590 7455 7642
rect 7455 7590 7501 7642
rect 7205 7588 7261 7590
rect 7285 7588 7341 7590
rect 7365 7588 7421 7590
rect 7445 7588 7501 7590
rect 7205 6554 7261 6556
rect 7285 6554 7341 6556
rect 7365 6554 7421 6556
rect 7445 6554 7501 6556
rect 7205 6502 7251 6554
rect 7251 6502 7261 6554
rect 7285 6502 7315 6554
rect 7315 6502 7327 6554
rect 7327 6502 7341 6554
rect 7365 6502 7379 6554
rect 7379 6502 7391 6554
rect 7391 6502 7421 6554
rect 7445 6502 7455 6554
rect 7455 6502 7501 6554
rect 7205 6500 7261 6502
rect 7285 6500 7341 6502
rect 7365 6500 7421 6502
rect 7445 6500 7501 6502
rect 6545 6010 6601 6012
rect 6625 6010 6681 6012
rect 6705 6010 6761 6012
rect 6785 6010 6841 6012
rect 6545 5958 6591 6010
rect 6591 5958 6601 6010
rect 6625 5958 6655 6010
rect 6655 5958 6667 6010
rect 6667 5958 6681 6010
rect 6705 5958 6719 6010
rect 6719 5958 6731 6010
rect 6731 5958 6761 6010
rect 6785 5958 6795 6010
rect 6795 5958 6841 6010
rect 6545 5956 6601 5958
rect 6625 5956 6681 5958
rect 6705 5956 6761 5958
rect 6785 5956 6841 5958
rect 6545 4922 6601 4924
rect 6625 4922 6681 4924
rect 6705 4922 6761 4924
rect 6785 4922 6841 4924
rect 6545 4870 6591 4922
rect 6591 4870 6601 4922
rect 6625 4870 6655 4922
rect 6655 4870 6667 4922
rect 6667 4870 6681 4922
rect 6705 4870 6719 4922
rect 6719 4870 6731 4922
rect 6731 4870 6761 4922
rect 6785 4870 6795 4922
rect 6795 4870 6841 4922
rect 6545 4868 6601 4870
rect 6625 4868 6681 4870
rect 6705 4868 6761 4870
rect 6785 4868 6841 4870
rect 7205 5466 7261 5468
rect 7285 5466 7341 5468
rect 7365 5466 7421 5468
rect 7445 5466 7501 5468
rect 7205 5414 7251 5466
rect 7251 5414 7261 5466
rect 7285 5414 7315 5466
rect 7315 5414 7327 5466
rect 7327 5414 7341 5466
rect 7365 5414 7379 5466
rect 7379 5414 7391 5466
rect 7391 5414 7421 5466
rect 7445 5414 7455 5466
rect 7455 5414 7501 5466
rect 7205 5412 7261 5414
rect 7285 5412 7341 5414
rect 7365 5412 7421 5414
rect 7445 5412 7501 5414
rect 6545 3834 6601 3836
rect 6625 3834 6681 3836
rect 6705 3834 6761 3836
rect 6785 3834 6841 3836
rect 6545 3782 6591 3834
rect 6591 3782 6601 3834
rect 6625 3782 6655 3834
rect 6655 3782 6667 3834
rect 6667 3782 6681 3834
rect 6705 3782 6719 3834
rect 6719 3782 6731 3834
rect 6731 3782 6761 3834
rect 6785 3782 6795 3834
rect 6795 3782 6841 3834
rect 6545 3780 6601 3782
rect 6625 3780 6681 3782
rect 6705 3780 6761 3782
rect 6785 3780 6841 3782
rect 7205 4378 7261 4380
rect 7285 4378 7341 4380
rect 7365 4378 7421 4380
rect 7445 4378 7501 4380
rect 7205 4326 7251 4378
rect 7251 4326 7261 4378
rect 7285 4326 7315 4378
rect 7315 4326 7327 4378
rect 7327 4326 7341 4378
rect 7365 4326 7379 4378
rect 7379 4326 7391 4378
rect 7391 4326 7421 4378
rect 7445 4326 7455 4378
rect 7455 4326 7501 4378
rect 7205 4324 7261 4326
rect 7285 4324 7341 4326
rect 7365 4324 7421 4326
rect 7445 4324 7501 4326
rect 7205 3290 7261 3292
rect 7285 3290 7341 3292
rect 7365 3290 7421 3292
rect 7445 3290 7501 3292
rect 7205 3238 7251 3290
rect 7251 3238 7261 3290
rect 7285 3238 7315 3290
rect 7315 3238 7327 3290
rect 7327 3238 7341 3290
rect 7365 3238 7379 3290
rect 7379 3238 7391 3290
rect 7391 3238 7421 3290
rect 7445 3238 7455 3290
rect 7455 3238 7501 3290
rect 7205 3236 7261 3238
rect 7285 3236 7341 3238
rect 7365 3236 7421 3238
rect 7445 3236 7501 3238
rect 10931 11994 10987 11996
rect 11011 11994 11067 11996
rect 11091 11994 11147 11996
rect 11171 11994 11227 11996
rect 10931 11942 10977 11994
rect 10977 11942 10987 11994
rect 11011 11942 11041 11994
rect 11041 11942 11053 11994
rect 11053 11942 11067 11994
rect 11091 11942 11105 11994
rect 11105 11942 11117 11994
rect 11117 11942 11147 11994
rect 11171 11942 11181 11994
rect 11181 11942 11227 11994
rect 10931 11940 10987 11942
rect 11011 11940 11067 11942
rect 11091 11940 11147 11942
rect 11171 11940 11227 11942
rect 14657 15258 14713 15260
rect 14737 15258 14793 15260
rect 14817 15258 14873 15260
rect 14897 15258 14953 15260
rect 14657 15206 14703 15258
rect 14703 15206 14713 15258
rect 14737 15206 14767 15258
rect 14767 15206 14779 15258
rect 14779 15206 14793 15258
rect 14817 15206 14831 15258
rect 14831 15206 14843 15258
rect 14843 15206 14873 15258
rect 14897 15206 14907 15258
rect 14907 15206 14953 15258
rect 14657 15204 14713 15206
rect 14737 15204 14793 15206
rect 14817 15204 14873 15206
rect 14897 15204 14953 15206
rect 13997 14714 14053 14716
rect 14077 14714 14133 14716
rect 14157 14714 14213 14716
rect 14237 14714 14293 14716
rect 13997 14662 14043 14714
rect 14043 14662 14053 14714
rect 14077 14662 14107 14714
rect 14107 14662 14119 14714
rect 14119 14662 14133 14714
rect 14157 14662 14171 14714
rect 14171 14662 14183 14714
rect 14183 14662 14213 14714
rect 14237 14662 14247 14714
rect 14247 14662 14293 14714
rect 13997 14660 14053 14662
rect 14077 14660 14133 14662
rect 14157 14660 14213 14662
rect 14237 14660 14293 14662
rect 14657 14170 14713 14172
rect 14737 14170 14793 14172
rect 14817 14170 14873 14172
rect 14897 14170 14953 14172
rect 14657 14118 14703 14170
rect 14703 14118 14713 14170
rect 14737 14118 14767 14170
rect 14767 14118 14779 14170
rect 14779 14118 14793 14170
rect 14817 14118 14831 14170
rect 14831 14118 14843 14170
rect 14843 14118 14873 14170
rect 14897 14118 14907 14170
rect 14907 14118 14953 14170
rect 14657 14116 14713 14118
rect 14737 14116 14793 14118
rect 14817 14116 14873 14118
rect 14897 14116 14953 14118
rect 13997 13626 14053 13628
rect 14077 13626 14133 13628
rect 14157 13626 14213 13628
rect 14237 13626 14293 13628
rect 13997 13574 14043 13626
rect 14043 13574 14053 13626
rect 14077 13574 14107 13626
rect 14107 13574 14119 13626
rect 14119 13574 14133 13626
rect 14157 13574 14171 13626
rect 14171 13574 14183 13626
rect 14183 13574 14213 13626
rect 14237 13574 14247 13626
rect 14247 13574 14293 13626
rect 13997 13572 14053 13574
rect 14077 13572 14133 13574
rect 14157 13572 14213 13574
rect 14237 13572 14293 13574
rect 10931 10906 10987 10908
rect 11011 10906 11067 10908
rect 11091 10906 11147 10908
rect 11171 10906 11227 10908
rect 10931 10854 10977 10906
rect 10977 10854 10987 10906
rect 11011 10854 11041 10906
rect 11041 10854 11053 10906
rect 11053 10854 11067 10906
rect 11091 10854 11105 10906
rect 11105 10854 11117 10906
rect 11117 10854 11147 10906
rect 11171 10854 11181 10906
rect 11181 10854 11227 10906
rect 10931 10852 10987 10854
rect 11011 10852 11067 10854
rect 11091 10852 11147 10854
rect 11171 10852 11227 10854
rect 10931 9818 10987 9820
rect 11011 9818 11067 9820
rect 11091 9818 11147 9820
rect 11171 9818 11227 9820
rect 10931 9766 10977 9818
rect 10977 9766 10987 9818
rect 11011 9766 11041 9818
rect 11041 9766 11053 9818
rect 11053 9766 11067 9818
rect 11091 9766 11105 9818
rect 11105 9766 11117 9818
rect 11117 9766 11147 9818
rect 11171 9766 11181 9818
rect 11181 9766 11227 9818
rect 10931 9764 10987 9766
rect 11011 9764 11067 9766
rect 11091 9764 11147 9766
rect 11171 9764 11227 9766
rect 10271 9274 10327 9276
rect 10351 9274 10407 9276
rect 10431 9274 10487 9276
rect 10511 9274 10567 9276
rect 10271 9222 10317 9274
rect 10317 9222 10327 9274
rect 10351 9222 10381 9274
rect 10381 9222 10393 9274
rect 10393 9222 10407 9274
rect 10431 9222 10445 9274
rect 10445 9222 10457 9274
rect 10457 9222 10487 9274
rect 10511 9222 10521 9274
rect 10521 9222 10567 9274
rect 10271 9220 10327 9222
rect 10351 9220 10407 9222
rect 10431 9220 10487 9222
rect 10511 9220 10567 9222
rect 10271 8186 10327 8188
rect 10351 8186 10407 8188
rect 10431 8186 10487 8188
rect 10511 8186 10567 8188
rect 10271 8134 10317 8186
rect 10317 8134 10327 8186
rect 10351 8134 10381 8186
rect 10381 8134 10393 8186
rect 10393 8134 10407 8186
rect 10431 8134 10445 8186
rect 10445 8134 10457 8186
rect 10457 8134 10487 8186
rect 10511 8134 10521 8186
rect 10521 8134 10567 8186
rect 10271 8132 10327 8134
rect 10351 8132 10407 8134
rect 10431 8132 10487 8134
rect 10511 8132 10567 8134
rect 10271 7098 10327 7100
rect 10351 7098 10407 7100
rect 10431 7098 10487 7100
rect 10511 7098 10567 7100
rect 10271 7046 10317 7098
rect 10317 7046 10327 7098
rect 10351 7046 10381 7098
rect 10381 7046 10393 7098
rect 10393 7046 10407 7098
rect 10431 7046 10445 7098
rect 10445 7046 10457 7098
rect 10457 7046 10487 7098
rect 10511 7046 10521 7098
rect 10521 7046 10567 7098
rect 10271 7044 10327 7046
rect 10351 7044 10407 7046
rect 10431 7044 10487 7046
rect 10511 7044 10567 7046
rect 10271 6010 10327 6012
rect 10351 6010 10407 6012
rect 10431 6010 10487 6012
rect 10511 6010 10567 6012
rect 10271 5958 10317 6010
rect 10317 5958 10327 6010
rect 10351 5958 10381 6010
rect 10381 5958 10393 6010
rect 10393 5958 10407 6010
rect 10431 5958 10445 6010
rect 10445 5958 10457 6010
rect 10457 5958 10487 6010
rect 10511 5958 10521 6010
rect 10521 5958 10567 6010
rect 10271 5956 10327 5958
rect 10351 5956 10407 5958
rect 10431 5956 10487 5958
rect 10511 5956 10567 5958
rect 11242 9036 11298 9072
rect 11242 9016 11244 9036
rect 11244 9016 11296 9036
rect 11296 9016 11298 9036
rect 11610 9052 11612 9072
rect 11612 9052 11664 9072
rect 11664 9052 11666 9072
rect 11610 9016 11666 9052
rect 10931 8730 10987 8732
rect 11011 8730 11067 8732
rect 11091 8730 11147 8732
rect 11171 8730 11227 8732
rect 10931 8678 10977 8730
rect 10977 8678 10987 8730
rect 11011 8678 11041 8730
rect 11041 8678 11053 8730
rect 11053 8678 11067 8730
rect 11091 8678 11105 8730
rect 11105 8678 11117 8730
rect 11117 8678 11147 8730
rect 11171 8678 11181 8730
rect 11181 8678 11227 8730
rect 10931 8676 10987 8678
rect 11011 8676 11067 8678
rect 11091 8676 11147 8678
rect 11171 8676 11227 8678
rect 10931 7642 10987 7644
rect 11011 7642 11067 7644
rect 11091 7642 11147 7644
rect 11171 7642 11227 7644
rect 10931 7590 10977 7642
rect 10977 7590 10987 7642
rect 11011 7590 11041 7642
rect 11041 7590 11053 7642
rect 11053 7590 11067 7642
rect 11091 7590 11105 7642
rect 11105 7590 11117 7642
rect 11117 7590 11147 7642
rect 11171 7590 11181 7642
rect 11181 7590 11227 7642
rect 10931 7588 10987 7590
rect 11011 7588 11067 7590
rect 11091 7588 11147 7590
rect 11171 7588 11227 7590
rect 10931 6554 10987 6556
rect 11011 6554 11067 6556
rect 11091 6554 11147 6556
rect 11171 6554 11227 6556
rect 10931 6502 10977 6554
rect 10977 6502 10987 6554
rect 11011 6502 11041 6554
rect 11041 6502 11053 6554
rect 11053 6502 11067 6554
rect 11091 6502 11105 6554
rect 11105 6502 11117 6554
rect 11117 6502 11147 6554
rect 11171 6502 11181 6554
rect 11181 6502 11227 6554
rect 10931 6500 10987 6502
rect 11011 6500 11067 6502
rect 11091 6500 11147 6502
rect 11171 6500 11227 6502
rect 10271 4922 10327 4924
rect 10351 4922 10407 4924
rect 10431 4922 10487 4924
rect 10511 4922 10567 4924
rect 10271 4870 10317 4922
rect 10317 4870 10327 4922
rect 10351 4870 10381 4922
rect 10381 4870 10393 4922
rect 10393 4870 10407 4922
rect 10431 4870 10445 4922
rect 10445 4870 10457 4922
rect 10457 4870 10487 4922
rect 10511 4870 10521 4922
rect 10521 4870 10567 4922
rect 10271 4868 10327 4870
rect 10351 4868 10407 4870
rect 10431 4868 10487 4870
rect 10511 4868 10567 4870
rect 10271 3834 10327 3836
rect 10351 3834 10407 3836
rect 10431 3834 10487 3836
rect 10511 3834 10567 3836
rect 10271 3782 10317 3834
rect 10317 3782 10327 3834
rect 10351 3782 10381 3834
rect 10381 3782 10393 3834
rect 10393 3782 10407 3834
rect 10431 3782 10445 3834
rect 10445 3782 10457 3834
rect 10457 3782 10487 3834
rect 10511 3782 10521 3834
rect 10521 3782 10567 3834
rect 10271 3780 10327 3782
rect 10351 3780 10407 3782
rect 10431 3780 10487 3782
rect 10511 3780 10567 3782
rect 13997 12538 14053 12540
rect 14077 12538 14133 12540
rect 14157 12538 14213 12540
rect 14237 12538 14293 12540
rect 13997 12486 14043 12538
rect 14043 12486 14053 12538
rect 14077 12486 14107 12538
rect 14107 12486 14119 12538
rect 14119 12486 14133 12538
rect 14157 12486 14171 12538
rect 14171 12486 14183 12538
rect 14183 12486 14213 12538
rect 14237 12486 14247 12538
rect 14247 12486 14293 12538
rect 13997 12484 14053 12486
rect 14077 12484 14133 12486
rect 14157 12484 14213 12486
rect 14237 12484 14293 12486
rect 14657 13082 14713 13084
rect 14737 13082 14793 13084
rect 14817 13082 14873 13084
rect 14897 13082 14953 13084
rect 14657 13030 14703 13082
rect 14703 13030 14713 13082
rect 14737 13030 14767 13082
rect 14767 13030 14779 13082
rect 14779 13030 14793 13082
rect 14817 13030 14831 13082
rect 14831 13030 14843 13082
rect 14843 13030 14873 13082
rect 14897 13030 14907 13082
rect 14907 13030 14953 13082
rect 14657 13028 14713 13030
rect 14737 13028 14793 13030
rect 14817 13028 14873 13030
rect 14897 13028 14953 13030
rect 13997 11450 14053 11452
rect 14077 11450 14133 11452
rect 14157 11450 14213 11452
rect 14237 11450 14293 11452
rect 13997 11398 14043 11450
rect 14043 11398 14053 11450
rect 14077 11398 14107 11450
rect 14107 11398 14119 11450
rect 14119 11398 14133 11450
rect 14157 11398 14171 11450
rect 14171 11398 14183 11450
rect 14183 11398 14213 11450
rect 14237 11398 14247 11450
rect 14247 11398 14293 11450
rect 13997 11396 14053 11398
rect 14077 11396 14133 11398
rect 14157 11396 14213 11398
rect 14237 11396 14293 11398
rect 14657 11994 14713 11996
rect 14737 11994 14793 11996
rect 14817 11994 14873 11996
rect 14897 11994 14953 11996
rect 14657 11942 14703 11994
rect 14703 11942 14713 11994
rect 14737 11942 14767 11994
rect 14767 11942 14779 11994
rect 14779 11942 14793 11994
rect 14817 11942 14831 11994
rect 14831 11942 14843 11994
rect 14843 11942 14873 11994
rect 14897 11942 14907 11994
rect 14907 11942 14953 11994
rect 14657 11940 14713 11942
rect 14737 11940 14793 11942
rect 14817 11940 14873 11942
rect 14897 11940 14953 11942
rect 13997 10362 14053 10364
rect 14077 10362 14133 10364
rect 14157 10362 14213 10364
rect 14237 10362 14293 10364
rect 13997 10310 14043 10362
rect 14043 10310 14053 10362
rect 14077 10310 14107 10362
rect 14107 10310 14119 10362
rect 14119 10310 14133 10362
rect 14157 10310 14171 10362
rect 14171 10310 14183 10362
rect 14183 10310 14213 10362
rect 14237 10310 14247 10362
rect 14247 10310 14293 10362
rect 13997 10308 14053 10310
rect 14077 10308 14133 10310
rect 14157 10308 14213 10310
rect 14237 10308 14293 10310
rect 14657 10906 14713 10908
rect 14737 10906 14793 10908
rect 14817 10906 14873 10908
rect 14897 10906 14953 10908
rect 14657 10854 14703 10906
rect 14703 10854 14713 10906
rect 14737 10854 14767 10906
rect 14767 10854 14779 10906
rect 14779 10854 14793 10906
rect 14817 10854 14831 10906
rect 14831 10854 14843 10906
rect 14843 10854 14873 10906
rect 14897 10854 14907 10906
rect 14907 10854 14953 10906
rect 14657 10852 14713 10854
rect 14737 10852 14793 10854
rect 14817 10852 14873 10854
rect 14897 10852 14953 10854
rect 13997 9274 14053 9276
rect 14077 9274 14133 9276
rect 14157 9274 14213 9276
rect 14237 9274 14293 9276
rect 13997 9222 14043 9274
rect 14043 9222 14053 9274
rect 14077 9222 14107 9274
rect 14107 9222 14119 9274
rect 14119 9222 14133 9274
rect 14157 9222 14171 9274
rect 14171 9222 14183 9274
rect 14183 9222 14213 9274
rect 14237 9222 14247 9274
rect 14247 9222 14293 9274
rect 13997 9220 14053 9222
rect 14077 9220 14133 9222
rect 14157 9220 14213 9222
rect 14237 9220 14293 9222
rect 13997 8186 14053 8188
rect 14077 8186 14133 8188
rect 14157 8186 14213 8188
rect 14237 8186 14293 8188
rect 13997 8134 14043 8186
rect 14043 8134 14053 8186
rect 14077 8134 14107 8186
rect 14107 8134 14119 8186
rect 14119 8134 14133 8186
rect 14157 8134 14171 8186
rect 14171 8134 14183 8186
rect 14183 8134 14213 8186
rect 14237 8134 14247 8186
rect 14247 8134 14293 8186
rect 13997 8132 14053 8134
rect 14077 8132 14133 8134
rect 14157 8132 14213 8134
rect 14237 8132 14293 8134
rect 10931 5466 10987 5468
rect 11011 5466 11067 5468
rect 11091 5466 11147 5468
rect 11171 5466 11227 5468
rect 10931 5414 10977 5466
rect 10977 5414 10987 5466
rect 11011 5414 11041 5466
rect 11041 5414 11053 5466
rect 11053 5414 11067 5466
rect 11091 5414 11105 5466
rect 11105 5414 11117 5466
rect 11117 5414 11147 5466
rect 11171 5414 11181 5466
rect 11181 5414 11227 5466
rect 10931 5412 10987 5414
rect 11011 5412 11067 5414
rect 11091 5412 11147 5414
rect 11171 5412 11227 5414
rect 10931 4378 10987 4380
rect 11011 4378 11067 4380
rect 11091 4378 11147 4380
rect 11171 4378 11227 4380
rect 10931 4326 10977 4378
rect 10977 4326 10987 4378
rect 11011 4326 11041 4378
rect 11041 4326 11053 4378
rect 11053 4326 11067 4378
rect 11091 4326 11105 4378
rect 11105 4326 11117 4378
rect 11117 4326 11147 4378
rect 11171 4326 11181 4378
rect 11181 4326 11227 4378
rect 10931 4324 10987 4326
rect 11011 4324 11067 4326
rect 11091 4324 11147 4326
rect 11171 4324 11227 4326
rect 10931 3290 10987 3292
rect 11011 3290 11067 3292
rect 11091 3290 11147 3292
rect 11171 3290 11227 3292
rect 10931 3238 10977 3290
rect 10977 3238 10987 3290
rect 11011 3238 11041 3290
rect 11041 3238 11053 3290
rect 11053 3238 11067 3290
rect 11091 3238 11105 3290
rect 11105 3238 11117 3290
rect 11117 3238 11147 3290
rect 11171 3238 11181 3290
rect 11181 3238 11227 3290
rect 10931 3236 10987 3238
rect 11011 3236 11067 3238
rect 11091 3236 11147 3238
rect 11171 3236 11227 3238
rect 14657 9818 14713 9820
rect 14737 9818 14793 9820
rect 14817 9818 14873 9820
rect 14897 9818 14953 9820
rect 14657 9766 14703 9818
rect 14703 9766 14713 9818
rect 14737 9766 14767 9818
rect 14767 9766 14779 9818
rect 14779 9766 14793 9818
rect 14817 9766 14831 9818
rect 14831 9766 14843 9818
rect 14843 9766 14873 9818
rect 14897 9766 14907 9818
rect 14907 9766 14953 9818
rect 14657 9764 14713 9766
rect 14737 9764 14793 9766
rect 14817 9764 14873 9766
rect 14897 9764 14953 9766
rect 13997 7098 14053 7100
rect 14077 7098 14133 7100
rect 14157 7098 14213 7100
rect 14237 7098 14293 7100
rect 13997 7046 14043 7098
rect 14043 7046 14053 7098
rect 14077 7046 14107 7098
rect 14107 7046 14119 7098
rect 14119 7046 14133 7098
rect 14157 7046 14171 7098
rect 14171 7046 14183 7098
rect 14183 7046 14213 7098
rect 14237 7046 14247 7098
rect 14247 7046 14293 7098
rect 13997 7044 14053 7046
rect 14077 7044 14133 7046
rect 14157 7044 14213 7046
rect 14237 7044 14293 7046
rect 13997 6010 14053 6012
rect 14077 6010 14133 6012
rect 14157 6010 14213 6012
rect 14237 6010 14293 6012
rect 13997 5958 14043 6010
rect 14043 5958 14053 6010
rect 14077 5958 14107 6010
rect 14107 5958 14119 6010
rect 14119 5958 14133 6010
rect 14157 5958 14171 6010
rect 14171 5958 14183 6010
rect 14183 5958 14213 6010
rect 14237 5958 14247 6010
rect 14247 5958 14293 6010
rect 13997 5956 14053 5958
rect 14077 5956 14133 5958
rect 14157 5956 14213 5958
rect 14237 5956 14293 5958
rect 13997 4922 14053 4924
rect 14077 4922 14133 4924
rect 14157 4922 14213 4924
rect 14237 4922 14293 4924
rect 13997 4870 14043 4922
rect 14043 4870 14053 4922
rect 14077 4870 14107 4922
rect 14107 4870 14119 4922
rect 14119 4870 14133 4922
rect 14157 4870 14171 4922
rect 14171 4870 14183 4922
rect 14183 4870 14213 4922
rect 14237 4870 14247 4922
rect 14247 4870 14293 4922
rect 13997 4868 14053 4870
rect 14077 4868 14133 4870
rect 14157 4868 14213 4870
rect 14237 4868 14293 4870
rect 14657 8730 14713 8732
rect 14737 8730 14793 8732
rect 14817 8730 14873 8732
rect 14897 8730 14953 8732
rect 14657 8678 14703 8730
rect 14703 8678 14713 8730
rect 14737 8678 14767 8730
rect 14767 8678 14779 8730
rect 14779 8678 14793 8730
rect 14817 8678 14831 8730
rect 14831 8678 14843 8730
rect 14843 8678 14873 8730
rect 14897 8678 14907 8730
rect 14907 8678 14953 8730
rect 14657 8676 14713 8678
rect 14737 8676 14793 8678
rect 14817 8676 14873 8678
rect 14897 8676 14953 8678
rect 14657 7642 14713 7644
rect 14737 7642 14793 7644
rect 14817 7642 14873 7644
rect 14897 7642 14953 7644
rect 14657 7590 14703 7642
rect 14703 7590 14713 7642
rect 14737 7590 14767 7642
rect 14767 7590 14779 7642
rect 14779 7590 14793 7642
rect 14817 7590 14831 7642
rect 14831 7590 14843 7642
rect 14843 7590 14873 7642
rect 14897 7590 14907 7642
rect 14907 7590 14953 7642
rect 14657 7588 14713 7590
rect 14737 7588 14793 7590
rect 14817 7588 14873 7590
rect 14897 7588 14953 7590
rect 16026 8900 16082 8936
rect 16026 8880 16028 8900
rect 16028 8880 16080 8900
rect 16080 8880 16082 8900
rect 14657 6554 14713 6556
rect 14737 6554 14793 6556
rect 14817 6554 14873 6556
rect 14897 6554 14953 6556
rect 14657 6502 14703 6554
rect 14703 6502 14713 6554
rect 14737 6502 14767 6554
rect 14767 6502 14779 6554
rect 14779 6502 14793 6554
rect 14817 6502 14831 6554
rect 14831 6502 14843 6554
rect 14843 6502 14873 6554
rect 14897 6502 14907 6554
rect 14907 6502 14953 6554
rect 14657 6500 14713 6502
rect 14737 6500 14793 6502
rect 14817 6500 14873 6502
rect 14897 6500 14953 6502
rect 14657 5466 14713 5468
rect 14737 5466 14793 5468
rect 14817 5466 14873 5468
rect 14897 5466 14953 5468
rect 14657 5414 14703 5466
rect 14703 5414 14713 5466
rect 14737 5414 14767 5466
rect 14767 5414 14779 5466
rect 14779 5414 14793 5466
rect 14817 5414 14831 5466
rect 14831 5414 14843 5466
rect 14843 5414 14873 5466
rect 14897 5414 14907 5466
rect 14907 5414 14953 5466
rect 14657 5412 14713 5414
rect 14737 5412 14793 5414
rect 14817 5412 14873 5414
rect 14897 5412 14953 5414
rect 2819 2746 2875 2748
rect 2899 2746 2955 2748
rect 2979 2746 3035 2748
rect 3059 2746 3115 2748
rect 2819 2694 2865 2746
rect 2865 2694 2875 2746
rect 2899 2694 2929 2746
rect 2929 2694 2941 2746
rect 2941 2694 2955 2746
rect 2979 2694 2993 2746
rect 2993 2694 3005 2746
rect 3005 2694 3035 2746
rect 3059 2694 3069 2746
rect 3069 2694 3115 2746
rect 2819 2692 2875 2694
rect 2899 2692 2955 2694
rect 2979 2692 3035 2694
rect 3059 2692 3115 2694
rect 6545 2746 6601 2748
rect 6625 2746 6681 2748
rect 6705 2746 6761 2748
rect 6785 2746 6841 2748
rect 6545 2694 6591 2746
rect 6591 2694 6601 2746
rect 6625 2694 6655 2746
rect 6655 2694 6667 2746
rect 6667 2694 6681 2746
rect 6705 2694 6719 2746
rect 6719 2694 6731 2746
rect 6731 2694 6761 2746
rect 6785 2694 6795 2746
rect 6795 2694 6841 2746
rect 6545 2692 6601 2694
rect 6625 2692 6681 2694
rect 6705 2692 6761 2694
rect 6785 2692 6841 2694
rect 10271 2746 10327 2748
rect 10351 2746 10407 2748
rect 10431 2746 10487 2748
rect 10511 2746 10567 2748
rect 10271 2694 10317 2746
rect 10317 2694 10327 2746
rect 10351 2694 10381 2746
rect 10381 2694 10393 2746
rect 10393 2694 10407 2746
rect 10431 2694 10445 2746
rect 10445 2694 10457 2746
rect 10457 2694 10487 2746
rect 10511 2694 10521 2746
rect 10521 2694 10567 2746
rect 10271 2692 10327 2694
rect 10351 2692 10407 2694
rect 10431 2692 10487 2694
rect 10511 2692 10567 2694
rect 14657 4378 14713 4380
rect 14737 4378 14793 4380
rect 14817 4378 14873 4380
rect 14897 4378 14953 4380
rect 14657 4326 14703 4378
rect 14703 4326 14713 4378
rect 14737 4326 14767 4378
rect 14767 4326 14779 4378
rect 14779 4326 14793 4378
rect 14817 4326 14831 4378
rect 14831 4326 14843 4378
rect 14843 4326 14873 4378
rect 14897 4326 14907 4378
rect 14907 4326 14953 4378
rect 14657 4324 14713 4326
rect 14737 4324 14793 4326
rect 14817 4324 14873 4326
rect 14897 4324 14953 4326
rect 13997 3834 14053 3836
rect 14077 3834 14133 3836
rect 14157 3834 14213 3836
rect 14237 3834 14293 3836
rect 13997 3782 14043 3834
rect 14043 3782 14053 3834
rect 14077 3782 14107 3834
rect 14107 3782 14119 3834
rect 14119 3782 14133 3834
rect 14157 3782 14171 3834
rect 14171 3782 14183 3834
rect 14183 3782 14213 3834
rect 14237 3782 14247 3834
rect 14247 3782 14293 3834
rect 13997 3780 14053 3782
rect 14077 3780 14133 3782
rect 14157 3780 14213 3782
rect 14237 3780 14293 3782
rect 14657 3290 14713 3292
rect 14737 3290 14793 3292
rect 14817 3290 14873 3292
rect 14897 3290 14953 3292
rect 14657 3238 14703 3290
rect 14703 3238 14713 3290
rect 14737 3238 14767 3290
rect 14767 3238 14779 3290
rect 14779 3238 14793 3290
rect 14817 3238 14831 3290
rect 14831 3238 14843 3290
rect 14843 3238 14873 3290
rect 14897 3238 14907 3290
rect 14907 3238 14953 3290
rect 14657 3236 14713 3238
rect 14737 3236 14793 3238
rect 14817 3236 14873 3238
rect 14897 3236 14953 3238
rect 13997 2746 14053 2748
rect 14077 2746 14133 2748
rect 14157 2746 14213 2748
rect 14237 2746 14293 2748
rect 13997 2694 14043 2746
rect 14043 2694 14053 2746
rect 14077 2694 14107 2746
rect 14107 2694 14119 2746
rect 14119 2694 14133 2746
rect 14157 2694 14171 2746
rect 14171 2694 14183 2746
rect 14183 2694 14213 2746
rect 14237 2694 14247 2746
rect 14247 2694 14293 2746
rect 13997 2692 14053 2694
rect 14077 2692 14133 2694
rect 14157 2692 14213 2694
rect 14237 2692 14293 2694
rect 3479 2202 3535 2204
rect 3559 2202 3615 2204
rect 3639 2202 3695 2204
rect 3719 2202 3775 2204
rect 3479 2150 3525 2202
rect 3525 2150 3535 2202
rect 3559 2150 3589 2202
rect 3589 2150 3601 2202
rect 3601 2150 3615 2202
rect 3639 2150 3653 2202
rect 3653 2150 3665 2202
rect 3665 2150 3695 2202
rect 3719 2150 3729 2202
rect 3729 2150 3775 2202
rect 3479 2148 3535 2150
rect 3559 2148 3615 2150
rect 3639 2148 3695 2150
rect 3719 2148 3775 2150
rect 7205 2202 7261 2204
rect 7285 2202 7341 2204
rect 7365 2202 7421 2204
rect 7445 2202 7501 2204
rect 7205 2150 7251 2202
rect 7251 2150 7261 2202
rect 7285 2150 7315 2202
rect 7315 2150 7327 2202
rect 7327 2150 7341 2202
rect 7365 2150 7379 2202
rect 7379 2150 7391 2202
rect 7391 2150 7421 2202
rect 7445 2150 7455 2202
rect 7455 2150 7501 2202
rect 7205 2148 7261 2150
rect 7285 2148 7341 2150
rect 7365 2148 7421 2150
rect 7445 2148 7501 2150
rect 10931 2202 10987 2204
rect 11011 2202 11067 2204
rect 11091 2202 11147 2204
rect 11171 2202 11227 2204
rect 10931 2150 10977 2202
rect 10977 2150 10987 2202
rect 11011 2150 11041 2202
rect 11041 2150 11053 2202
rect 11053 2150 11067 2202
rect 11091 2150 11105 2202
rect 11105 2150 11117 2202
rect 11117 2150 11147 2202
rect 11171 2150 11181 2202
rect 11181 2150 11227 2202
rect 10931 2148 10987 2150
rect 11011 2148 11067 2150
rect 11091 2148 11147 2150
rect 11171 2148 11227 2150
rect 14657 2202 14713 2204
rect 14737 2202 14793 2204
rect 14817 2202 14873 2204
rect 14897 2202 14953 2204
rect 14657 2150 14703 2202
rect 14703 2150 14713 2202
rect 14737 2150 14767 2202
rect 14767 2150 14779 2202
rect 14779 2150 14793 2202
rect 14817 2150 14831 2202
rect 14831 2150 14843 2202
rect 14843 2150 14873 2202
rect 14897 2150 14907 2202
rect 14907 2150 14953 2202
rect 14657 2148 14713 2150
rect 14737 2148 14793 2150
rect 14817 2148 14873 2150
rect 14897 2148 14953 2150
<< metal3 >>
rect 0 17008 800 17128
rect 2809 16896 3125 16897
rect 2809 16832 2815 16896
rect 2879 16832 2895 16896
rect 2959 16832 2975 16896
rect 3039 16832 3055 16896
rect 3119 16832 3125 16896
rect 2809 16831 3125 16832
rect 6535 16896 6851 16897
rect 6535 16832 6541 16896
rect 6605 16832 6621 16896
rect 6685 16832 6701 16896
rect 6765 16832 6781 16896
rect 6845 16832 6851 16896
rect 6535 16831 6851 16832
rect 10261 16896 10577 16897
rect 10261 16832 10267 16896
rect 10331 16832 10347 16896
rect 10411 16832 10427 16896
rect 10491 16832 10507 16896
rect 10571 16832 10577 16896
rect 10261 16831 10577 16832
rect 13987 16896 14303 16897
rect 13987 16832 13993 16896
rect 14057 16832 14073 16896
rect 14137 16832 14153 16896
rect 14217 16832 14233 16896
rect 14297 16832 14303 16896
rect 13987 16831 14303 16832
rect 3469 16352 3785 16353
rect 3469 16288 3475 16352
rect 3539 16288 3555 16352
rect 3619 16288 3635 16352
rect 3699 16288 3715 16352
rect 3779 16288 3785 16352
rect 3469 16287 3785 16288
rect 7195 16352 7511 16353
rect 7195 16288 7201 16352
rect 7265 16288 7281 16352
rect 7345 16288 7361 16352
rect 7425 16288 7441 16352
rect 7505 16288 7511 16352
rect 7195 16287 7511 16288
rect 10921 16352 11237 16353
rect 10921 16288 10927 16352
rect 10991 16288 11007 16352
rect 11071 16288 11087 16352
rect 11151 16288 11167 16352
rect 11231 16288 11237 16352
rect 10921 16287 11237 16288
rect 14647 16352 14963 16353
rect 14647 16288 14653 16352
rect 14717 16288 14733 16352
rect 14797 16288 14813 16352
rect 14877 16288 14893 16352
rect 14957 16288 14963 16352
rect 14647 16287 14963 16288
rect 2809 15808 3125 15809
rect 2809 15744 2815 15808
rect 2879 15744 2895 15808
rect 2959 15744 2975 15808
rect 3039 15744 3055 15808
rect 3119 15744 3125 15808
rect 2809 15743 3125 15744
rect 6535 15808 6851 15809
rect 6535 15744 6541 15808
rect 6605 15744 6621 15808
rect 6685 15744 6701 15808
rect 6765 15744 6781 15808
rect 6845 15744 6851 15808
rect 6535 15743 6851 15744
rect 10261 15808 10577 15809
rect 10261 15744 10267 15808
rect 10331 15744 10347 15808
rect 10411 15744 10427 15808
rect 10491 15744 10507 15808
rect 10571 15744 10577 15808
rect 10261 15743 10577 15744
rect 13987 15808 14303 15809
rect 13987 15744 13993 15808
rect 14057 15744 14073 15808
rect 14137 15744 14153 15808
rect 14217 15744 14233 15808
rect 14297 15744 14303 15808
rect 13987 15743 14303 15744
rect 16402 15648 17202 15768
rect 3469 15264 3785 15265
rect 3469 15200 3475 15264
rect 3539 15200 3555 15264
rect 3619 15200 3635 15264
rect 3699 15200 3715 15264
rect 3779 15200 3785 15264
rect 3469 15199 3785 15200
rect 7195 15264 7511 15265
rect 7195 15200 7201 15264
rect 7265 15200 7281 15264
rect 7345 15200 7361 15264
rect 7425 15200 7441 15264
rect 7505 15200 7511 15264
rect 7195 15199 7511 15200
rect 10921 15264 11237 15265
rect 10921 15200 10927 15264
rect 10991 15200 11007 15264
rect 11071 15200 11087 15264
rect 11151 15200 11167 15264
rect 11231 15200 11237 15264
rect 10921 15199 11237 15200
rect 14647 15264 14963 15265
rect 14647 15200 14653 15264
rect 14717 15200 14733 15264
rect 14797 15200 14813 15264
rect 14877 15200 14893 15264
rect 14957 15200 14963 15264
rect 14647 15199 14963 15200
rect 2809 14720 3125 14721
rect 2809 14656 2815 14720
rect 2879 14656 2895 14720
rect 2959 14656 2975 14720
rect 3039 14656 3055 14720
rect 3119 14656 3125 14720
rect 2809 14655 3125 14656
rect 6535 14720 6851 14721
rect 6535 14656 6541 14720
rect 6605 14656 6621 14720
rect 6685 14656 6701 14720
rect 6765 14656 6781 14720
rect 6845 14656 6851 14720
rect 6535 14655 6851 14656
rect 10261 14720 10577 14721
rect 10261 14656 10267 14720
rect 10331 14656 10347 14720
rect 10411 14656 10427 14720
rect 10491 14656 10507 14720
rect 10571 14656 10577 14720
rect 10261 14655 10577 14656
rect 13987 14720 14303 14721
rect 13987 14656 13993 14720
rect 14057 14656 14073 14720
rect 14137 14656 14153 14720
rect 14217 14656 14233 14720
rect 14297 14656 14303 14720
rect 13987 14655 14303 14656
rect 3469 14176 3785 14177
rect 3469 14112 3475 14176
rect 3539 14112 3555 14176
rect 3619 14112 3635 14176
rect 3699 14112 3715 14176
rect 3779 14112 3785 14176
rect 3469 14111 3785 14112
rect 7195 14176 7511 14177
rect 7195 14112 7201 14176
rect 7265 14112 7281 14176
rect 7345 14112 7361 14176
rect 7425 14112 7441 14176
rect 7505 14112 7511 14176
rect 7195 14111 7511 14112
rect 10921 14176 11237 14177
rect 10921 14112 10927 14176
rect 10991 14112 11007 14176
rect 11071 14112 11087 14176
rect 11151 14112 11167 14176
rect 11231 14112 11237 14176
rect 10921 14111 11237 14112
rect 14647 14176 14963 14177
rect 14647 14112 14653 14176
rect 14717 14112 14733 14176
rect 14797 14112 14813 14176
rect 14877 14112 14893 14176
rect 14957 14112 14963 14176
rect 14647 14111 14963 14112
rect 0 13608 800 13728
rect 2809 13632 3125 13633
rect 2809 13568 2815 13632
rect 2879 13568 2895 13632
rect 2959 13568 2975 13632
rect 3039 13568 3055 13632
rect 3119 13568 3125 13632
rect 2809 13567 3125 13568
rect 6535 13632 6851 13633
rect 6535 13568 6541 13632
rect 6605 13568 6621 13632
rect 6685 13568 6701 13632
rect 6765 13568 6781 13632
rect 6845 13568 6851 13632
rect 6535 13567 6851 13568
rect 10261 13632 10577 13633
rect 10261 13568 10267 13632
rect 10331 13568 10347 13632
rect 10411 13568 10427 13632
rect 10491 13568 10507 13632
rect 10571 13568 10577 13632
rect 10261 13567 10577 13568
rect 13987 13632 14303 13633
rect 13987 13568 13993 13632
rect 14057 13568 14073 13632
rect 14137 13568 14153 13632
rect 14217 13568 14233 13632
rect 14297 13568 14303 13632
rect 13987 13567 14303 13568
rect 3469 13088 3785 13089
rect 3469 13024 3475 13088
rect 3539 13024 3555 13088
rect 3619 13024 3635 13088
rect 3699 13024 3715 13088
rect 3779 13024 3785 13088
rect 3469 13023 3785 13024
rect 7195 13088 7511 13089
rect 7195 13024 7201 13088
rect 7265 13024 7281 13088
rect 7345 13024 7361 13088
rect 7425 13024 7441 13088
rect 7505 13024 7511 13088
rect 7195 13023 7511 13024
rect 10921 13088 11237 13089
rect 10921 13024 10927 13088
rect 10991 13024 11007 13088
rect 11071 13024 11087 13088
rect 11151 13024 11167 13088
rect 11231 13024 11237 13088
rect 10921 13023 11237 13024
rect 14647 13088 14963 13089
rect 14647 13024 14653 13088
rect 14717 13024 14733 13088
rect 14797 13024 14813 13088
rect 14877 13024 14893 13088
rect 14957 13024 14963 13088
rect 14647 13023 14963 13024
rect 2809 12544 3125 12545
rect 2809 12480 2815 12544
rect 2879 12480 2895 12544
rect 2959 12480 2975 12544
rect 3039 12480 3055 12544
rect 3119 12480 3125 12544
rect 2809 12479 3125 12480
rect 6535 12544 6851 12545
rect 6535 12480 6541 12544
rect 6605 12480 6621 12544
rect 6685 12480 6701 12544
rect 6765 12480 6781 12544
rect 6845 12480 6851 12544
rect 6535 12479 6851 12480
rect 10261 12544 10577 12545
rect 10261 12480 10267 12544
rect 10331 12480 10347 12544
rect 10411 12480 10427 12544
rect 10491 12480 10507 12544
rect 10571 12480 10577 12544
rect 10261 12479 10577 12480
rect 13987 12544 14303 12545
rect 13987 12480 13993 12544
rect 14057 12480 14073 12544
rect 14137 12480 14153 12544
rect 14217 12480 14233 12544
rect 14297 12480 14303 12544
rect 13987 12479 14303 12480
rect 16402 12248 17202 12368
rect 3469 12000 3785 12001
rect 3469 11936 3475 12000
rect 3539 11936 3555 12000
rect 3619 11936 3635 12000
rect 3699 11936 3715 12000
rect 3779 11936 3785 12000
rect 3469 11935 3785 11936
rect 7195 12000 7511 12001
rect 7195 11936 7201 12000
rect 7265 11936 7281 12000
rect 7345 11936 7361 12000
rect 7425 11936 7441 12000
rect 7505 11936 7511 12000
rect 7195 11935 7511 11936
rect 10921 12000 11237 12001
rect 10921 11936 10927 12000
rect 10991 11936 11007 12000
rect 11071 11936 11087 12000
rect 11151 11936 11167 12000
rect 11231 11936 11237 12000
rect 10921 11935 11237 11936
rect 14647 12000 14963 12001
rect 14647 11936 14653 12000
rect 14717 11936 14733 12000
rect 14797 11936 14813 12000
rect 14877 11936 14893 12000
rect 14957 11936 14963 12000
rect 14647 11935 14963 11936
rect 2809 11456 3125 11457
rect 2809 11392 2815 11456
rect 2879 11392 2895 11456
rect 2959 11392 2975 11456
rect 3039 11392 3055 11456
rect 3119 11392 3125 11456
rect 2809 11391 3125 11392
rect 6535 11456 6851 11457
rect 6535 11392 6541 11456
rect 6605 11392 6621 11456
rect 6685 11392 6701 11456
rect 6765 11392 6781 11456
rect 6845 11392 6851 11456
rect 6535 11391 6851 11392
rect 10261 11456 10577 11457
rect 10261 11392 10267 11456
rect 10331 11392 10347 11456
rect 10411 11392 10427 11456
rect 10491 11392 10507 11456
rect 10571 11392 10577 11456
rect 10261 11391 10577 11392
rect 13987 11456 14303 11457
rect 13987 11392 13993 11456
rect 14057 11392 14073 11456
rect 14137 11392 14153 11456
rect 14217 11392 14233 11456
rect 14297 11392 14303 11456
rect 13987 11391 14303 11392
rect 3469 10912 3785 10913
rect 3469 10848 3475 10912
rect 3539 10848 3555 10912
rect 3619 10848 3635 10912
rect 3699 10848 3715 10912
rect 3779 10848 3785 10912
rect 3469 10847 3785 10848
rect 7195 10912 7511 10913
rect 7195 10848 7201 10912
rect 7265 10848 7281 10912
rect 7345 10848 7361 10912
rect 7425 10848 7441 10912
rect 7505 10848 7511 10912
rect 7195 10847 7511 10848
rect 10921 10912 11237 10913
rect 10921 10848 10927 10912
rect 10991 10848 11007 10912
rect 11071 10848 11087 10912
rect 11151 10848 11167 10912
rect 11231 10848 11237 10912
rect 10921 10847 11237 10848
rect 14647 10912 14963 10913
rect 14647 10848 14653 10912
rect 14717 10848 14733 10912
rect 14797 10848 14813 10912
rect 14877 10848 14893 10912
rect 14957 10848 14963 10912
rect 14647 10847 14963 10848
rect 2809 10368 3125 10369
rect 0 10298 800 10328
rect 2809 10304 2815 10368
rect 2879 10304 2895 10368
rect 2959 10304 2975 10368
rect 3039 10304 3055 10368
rect 3119 10304 3125 10368
rect 2809 10303 3125 10304
rect 6535 10368 6851 10369
rect 6535 10304 6541 10368
rect 6605 10304 6621 10368
rect 6685 10304 6701 10368
rect 6765 10304 6781 10368
rect 6845 10304 6851 10368
rect 6535 10303 6851 10304
rect 10261 10368 10577 10369
rect 10261 10304 10267 10368
rect 10331 10304 10347 10368
rect 10411 10304 10427 10368
rect 10491 10304 10507 10368
rect 10571 10304 10577 10368
rect 10261 10303 10577 10304
rect 13987 10368 14303 10369
rect 13987 10304 13993 10368
rect 14057 10304 14073 10368
rect 14137 10304 14153 10368
rect 14217 10304 14233 10368
rect 14297 10304 14303 10368
rect 13987 10303 14303 10304
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10208 800 10238
rect 933 10235 999 10238
rect 3469 9824 3785 9825
rect 3469 9760 3475 9824
rect 3539 9760 3555 9824
rect 3619 9760 3635 9824
rect 3699 9760 3715 9824
rect 3779 9760 3785 9824
rect 3469 9759 3785 9760
rect 7195 9824 7511 9825
rect 7195 9760 7201 9824
rect 7265 9760 7281 9824
rect 7345 9760 7361 9824
rect 7425 9760 7441 9824
rect 7505 9760 7511 9824
rect 7195 9759 7511 9760
rect 10921 9824 11237 9825
rect 10921 9760 10927 9824
rect 10991 9760 11007 9824
rect 11071 9760 11087 9824
rect 11151 9760 11167 9824
rect 11231 9760 11237 9824
rect 10921 9759 11237 9760
rect 14647 9824 14963 9825
rect 14647 9760 14653 9824
rect 14717 9760 14733 9824
rect 14797 9760 14813 9824
rect 14877 9760 14893 9824
rect 14957 9760 14963 9824
rect 14647 9759 14963 9760
rect 657 9618 723 9621
rect 8753 9618 8819 9621
rect 657 9616 8819 9618
rect 657 9560 662 9616
rect 718 9560 8758 9616
rect 8814 9560 8819 9616
rect 657 9558 8819 9560
rect 657 9555 723 9558
rect 8753 9555 8819 9558
rect 2809 9280 3125 9281
rect 2809 9216 2815 9280
rect 2879 9216 2895 9280
rect 2959 9216 2975 9280
rect 3039 9216 3055 9280
rect 3119 9216 3125 9280
rect 2809 9215 3125 9216
rect 6535 9280 6851 9281
rect 6535 9216 6541 9280
rect 6605 9216 6621 9280
rect 6685 9216 6701 9280
rect 6765 9216 6781 9280
rect 6845 9216 6851 9280
rect 6535 9215 6851 9216
rect 10261 9280 10577 9281
rect 10261 9216 10267 9280
rect 10331 9216 10347 9280
rect 10411 9216 10427 9280
rect 10491 9216 10507 9280
rect 10571 9216 10577 9280
rect 10261 9215 10577 9216
rect 13987 9280 14303 9281
rect 13987 9216 13993 9280
rect 14057 9216 14073 9280
rect 14137 9216 14153 9280
rect 14217 9216 14233 9280
rect 14297 9216 14303 9280
rect 13987 9215 14303 9216
rect 11237 9074 11303 9077
rect 11605 9074 11671 9077
rect 11237 9072 11671 9074
rect 11237 9016 11242 9072
rect 11298 9016 11610 9072
rect 11666 9016 11671 9072
rect 11237 9014 11671 9016
rect 11237 9011 11303 9014
rect 11605 9011 11671 9014
rect 16021 8938 16087 8941
rect 16402 8938 17202 8968
rect 16021 8936 17202 8938
rect 16021 8880 16026 8936
rect 16082 8880 17202 8936
rect 16021 8878 17202 8880
rect 16021 8875 16087 8878
rect 16402 8848 17202 8878
rect 3469 8736 3785 8737
rect 3469 8672 3475 8736
rect 3539 8672 3555 8736
rect 3619 8672 3635 8736
rect 3699 8672 3715 8736
rect 3779 8672 3785 8736
rect 3469 8671 3785 8672
rect 7195 8736 7511 8737
rect 7195 8672 7201 8736
rect 7265 8672 7281 8736
rect 7345 8672 7361 8736
rect 7425 8672 7441 8736
rect 7505 8672 7511 8736
rect 7195 8671 7511 8672
rect 10921 8736 11237 8737
rect 10921 8672 10927 8736
rect 10991 8672 11007 8736
rect 11071 8672 11087 8736
rect 11151 8672 11167 8736
rect 11231 8672 11237 8736
rect 10921 8671 11237 8672
rect 14647 8736 14963 8737
rect 14647 8672 14653 8736
rect 14717 8672 14733 8736
rect 14797 8672 14813 8736
rect 14877 8672 14893 8736
rect 14957 8672 14963 8736
rect 14647 8671 14963 8672
rect 2809 8192 3125 8193
rect 2809 8128 2815 8192
rect 2879 8128 2895 8192
rect 2959 8128 2975 8192
rect 3039 8128 3055 8192
rect 3119 8128 3125 8192
rect 2809 8127 3125 8128
rect 6535 8192 6851 8193
rect 6535 8128 6541 8192
rect 6605 8128 6621 8192
rect 6685 8128 6701 8192
rect 6765 8128 6781 8192
rect 6845 8128 6851 8192
rect 6535 8127 6851 8128
rect 10261 8192 10577 8193
rect 10261 8128 10267 8192
rect 10331 8128 10347 8192
rect 10411 8128 10427 8192
rect 10491 8128 10507 8192
rect 10571 8128 10577 8192
rect 10261 8127 10577 8128
rect 13987 8192 14303 8193
rect 13987 8128 13993 8192
rect 14057 8128 14073 8192
rect 14137 8128 14153 8192
rect 14217 8128 14233 8192
rect 14297 8128 14303 8192
rect 13987 8127 14303 8128
rect 3469 7648 3785 7649
rect 3469 7584 3475 7648
rect 3539 7584 3555 7648
rect 3619 7584 3635 7648
rect 3699 7584 3715 7648
rect 3779 7584 3785 7648
rect 3469 7583 3785 7584
rect 7195 7648 7511 7649
rect 7195 7584 7201 7648
rect 7265 7584 7281 7648
rect 7345 7584 7361 7648
rect 7425 7584 7441 7648
rect 7505 7584 7511 7648
rect 7195 7583 7511 7584
rect 10921 7648 11237 7649
rect 10921 7584 10927 7648
rect 10991 7584 11007 7648
rect 11071 7584 11087 7648
rect 11151 7584 11167 7648
rect 11231 7584 11237 7648
rect 10921 7583 11237 7584
rect 14647 7648 14963 7649
rect 14647 7584 14653 7648
rect 14717 7584 14733 7648
rect 14797 7584 14813 7648
rect 14877 7584 14893 7648
rect 14957 7584 14963 7648
rect 14647 7583 14963 7584
rect 2809 7104 3125 7105
rect 2809 7040 2815 7104
rect 2879 7040 2895 7104
rect 2959 7040 2975 7104
rect 3039 7040 3055 7104
rect 3119 7040 3125 7104
rect 2809 7039 3125 7040
rect 6535 7104 6851 7105
rect 6535 7040 6541 7104
rect 6605 7040 6621 7104
rect 6685 7040 6701 7104
rect 6765 7040 6781 7104
rect 6845 7040 6851 7104
rect 6535 7039 6851 7040
rect 10261 7104 10577 7105
rect 10261 7040 10267 7104
rect 10331 7040 10347 7104
rect 10411 7040 10427 7104
rect 10491 7040 10507 7104
rect 10571 7040 10577 7104
rect 10261 7039 10577 7040
rect 13987 7104 14303 7105
rect 13987 7040 13993 7104
rect 14057 7040 14073 7104
rect 14137 7040 14153 7104
rect 14217 7040 14233 7104
rect 14297 7040 14303 7104
rect 13987 7039 14303 7040
rect 0 6808 800 6928
rect 3469 6560 3785 6561
rect 3469 6496 3475 6560
rect 3539 6496 3555 6560
rect 3619 6496 3635 6560
rect 3699 6496 3715 6560
rect 3779 6496 3785 6560
rect 3469 6495 3785 6496
rect 7195 6560 7511 6561
rect 7195 6496 7201 6560
rect 7265 6496 7281 6560
rect 7345 6496 7361 6560
rect 7425 6496 7441 6560
rect 7505 6496 7511 6560
rect 7195 6495 7511 6496
rect 10921 6560 11237 6561
rect 10921 6496 10927 6560
rect 10991 6496 11007 6560
rect 11071 6496 11087 6560
rect 11151 6496 11167 6560
rect 11231 6496 11237 6560
rect 10921 6495 11237 6496
rect 14647 6560 14963 6561
rect 14647 6496 14653 6560
rect 14717 6496 14733 6560
rect 14797 6496 14813 6560
rect 14877 6496 14893 6560
rect 14957 6496 14963 6560
rect 14647 6495 14963 6496
rect 2809 6016 3125 6017
rect 2809 5952 2815 6016
rect 2879 5952 2895 6016
rect 2959 5952 2975 6016
rect 3039 5952 3055 6016
rect 3119 5952 3125 6016
rect 2809 5951 3125 5952
rect 6535 6016 6851 6017
rect 6535 5952 6541 6016
rect 6605 5952 6621 6016
rect 6685 5952 6701 6016
rect 6765 5952 6781 6016
rect 6845 5952 6851 6016
rect 6535 5951 6851 5952
rect 10261 6016 10577 6017
rect 10261 5952 10267 6016
rect 10331 5952 10347 6016
rect 10411 5952 10427 6016
rect 10491 5952 10507 6016
rect 10571 5952 10577 6016
rect 10261 5951 10577 5952
rect 13987 6016 14303 6017
rect 13987 5952 13993 6016
rect 14057 5952 14073 6016
rect 14137 5952 14153 6016
rect 14217 5952 14233 6016
rect 14297 5952 14303 6016
rect 13987 5951 14303 5952
rect 3469 5472 3785 5473
rect 3469 5408 3475 5472
rect 3539 5408 3555 5472
rect 3619 5408 3635 5472
rect 3699 5408 3715 5472
rect 3779 5408 3785 5472
rect 3469 5407 3785 5408
rect 7195 5472 7511 5473
rect 7195 5408 7201 5472
rect 7265 5408 7281 5472
rect 7345 5408 7361 5472
rect 7425 5408 7441 5472
rect 7505 5408 7511 5472
rect 7195 5407 7511 5408
rect 10921 5472 11237 5473
rect 10921 5408 10927 5472
rect 10991 5408 11007 5472
rect 11071 5408 11087 5472
rect 11151 5408 11167 5472
rect 11231 5408 11237 5472
rect 10921 5407 11237 5408
rect 14647 5472 14963 5473
rect 14647 5408 14653 5472
rect 14717 5408 14733 5472
rect 14797 5408 14813 5472
rect 14877 5408 14893 5472
rect 14957 5408 14963 5472
rect 16402 5448 17202 5568
rect 14647 5407 14963 5408
rect 2809 4928 3125 4929
rect 2809 4864 2815 4928
rect 2879 4864 2895 4928
rect 2959 4864 2975 4928
rect 3039 4864 3055 4928
rect 3119 4864 3125 4928
rect 2809 4863 3125 4864
rect 6535 4928 6851 4929
rect 6535 4864 6541 4928
rect 6605 4864 6621 4928
rect 6685 4864 6701 4928
rect 6765 4864 6781 4928
rect 6845 4864 6851 4928
rect 6535 4863 6851 4864
rect 10261 4928 10577 4929
rect 10261 4864 10267 4928
rect 10331 4864 10347 4928
rect 10411 4864 10427 4928
rect 10491 4864 10507 4928
rect 10571 4864 10577 4928
rect 10261 4863 10577 4864
rect 13987 4928 14303 4929
rect 13987 4864 13993 4928
rect 14057 4864 14073 4928
rect 14137 4864 14153 4928
rect 14217 4864 14233 4928
rect 14297 4864 14303 4928
rect 13987 4863 14303 4864
rect 3469 4384 3785 4385
rect 3469 4320 3475 4384
rect 3539 4320 3555 4384
rect 3619 4320 3635 4384
rect 3699 4320 3715 4384
rect 3779 4320 3785 4384
rect 3469 4319 3785 4320
rect 7195 4384 7511 4385
rect 7195 4320 7201 4384
rect 7265 4320 7281 4384
rect 7345 4320 7361 4384
rect 7425 4320 7441 4384
rect 7505 4320 7511 4384
rect 7195 4319 7511 4320
rect 10921 4384 11237 4385
rect 10921 4320 10927 4384
rect 10991 4320 11007 4384
rect 11071 4320 11087 4384
rect 11151 4320 11167 4384
rect 11231 4320 11237 4384
rect 10921 4319 11237 4320
rect 14647 4384 14963 4385
rect 14647 4320 14653 4384
rect 14717 4320 14733 4384
rect 14797 4320 14813 4384
rect 14877 4320 14893 4384
rect 14957 4320 14963 4384
rect 14647 4319 14963 4320
rect 2809 3840 3125 3841
rect 2809 3776 2815 3840
rect 2879 3776 2895 3840
rect 2959 3776 2975 3840
rect 3039 3776 3055 3840
rect 3119 3776 3125 3840
rect 2809 3775 3125 3776
rect 6535 3840 6851 3841
rect 6535 3776 6541 3840
rect 6605 3776 6621 3840
rect 6685 3776 6701 3840
rect 6765 3776 6781 3840
rect 6845 3776 6851 3840
rect 6535 3775 6851 3776
rect 10261 3840 10577 3841
rect 10261 3776 10267 3840
rect 10331 3776 10347 3840
rect 10411 3776 10427 3840
rect 10491 3776 10507 3840
rect 10571 3776 10577 3840
rect 10261 3775 10577 3776
rect 13987 3840 14303 3841
rect 13987 3776 13993 3840
rect 14057 3776 14073 3840
rect 14137 3776 14153 3840
rect 14217 3776 14233 3840
rect 14297 3776 14303 3840
rect 13987 3775 14303 3776
rect 0 3408 800 3528
rect 3469 3296 3785 3297
rect 3469 3232 3475 3296
rect 3539 3232 3555 3296
rect 3619 3232 3635 3296
rect 3699 3232 3715 3296
rect 3779 3232 3785 3296
rect 3469 3231 3785 3232
rect 7195 3296 7511 3297
rect 7195 3232 7201 3296
rect 7265 3232 7281 3296
rect 7345 3232 7361 3296
rect 7425 3232 7441 3296
rect 7505 3232 7511 3296
rect 7195 3231 7511 3232
rect 10921 3296 11237 3297
rect 10921 3232 10927 3296
rect 10991 3232 11007 3296
rect 11071 3232 11087 3296
rect 11151 3232 11167 3296
rect 11231 3232 11237 3296
rect 10921 3231 11237 3232
rect 14647 3296 14963 3297
rect 14647 3232 14653 3296
rect 14717 3232 14733 3296
rect 14797 3232 14813 3296
rect 14877 3232 14893 3296
rect 14957 3232 14963 3296
rect 14647 3231 14963 3232
rect 2809 2752 3125 2753
rect 2809 2688 2815 2752
rect 2879 2688 2895 2752
rect 2959 2688 2975 2752
rect 3039 2688 3055 2752
rect 3119 2688 3125 2752
rect 2809 2687 3125 2688
rect 6535 2752 6851 2753
rect 6535 2688 6541 2752
rect 6605 2688 6621 2752
rect 6685 2688 6701 2752
rect 6765 2688 6781 2752
rect 6845 2688 6851 2752
rect 6535 2687 6851 2688
rect 10261 2752 10577 2753
rect 10261 2688 10267 2752
rect 10331 2688 10347 2752
rect 10411 2688 10427 2752
rect 10491 2688 10507 2752
rect 10571 2688 10577 2752
rect 10261 2687 10577 2688
rect 13987 2752 14303 2753
rect 13987 2688 13993 2752
rect 14057 2688 14073 2752
rect 14137 2688 14153 2752
rect 14217 2688 14233 2752
rect 14297 2688 14303 2752
rect 13987 2687 14303 2688
rect 3469 2208 3785 2209
rect 3469 2144 3475 2208
rect 3539 2144 3555 2208
rect 3619 2144 3635 2208
rect 3699 2144 3715 2208
rect 3779 2144 3785 2208
rect 3469 2143 3785 2144
rect 7195 2208 7511 2209
rect 7195 2144 7201 2208
rect 7265 2144 7281 2208
rect 7345 2144 7361 2208
rect 7425 2144 7441 2208
rect 7505 2144 7511 2208
rect 7195 2143 7511 2144
rect 10921 2208 11237 2209
rect 10921 2144 10927 2208
rect 10991 2144 11007 2208
rect 11071 2144 11087 2208
rect 11151 2144 11167 2208
rect 11231 2144 11237 2208
rect 10921 2143 11237 2144
rect 14647 2208 14963 2209
rect 14647 2144 14653 2208
rect 14717 2144 14733 2208
rect 14797 2144 14813 2208
rect 14877 2144 14893 2208
rect 14957 2144 14963 2208
rect 14647 2143 14963 2144
rect 16402 2048 17202 2168
<< via3 >>
rect 2815 16892 2879 16896
rect 2815 16836 2819 16892
rect 2819 16836 2875 16892
rect 2875 16836 2879 16892
rect 2815 16832 2879 16836
rect 2895 16892 2959 16896
rect 2895 16836 2899 16892
rect 2899 16836 2955 16892
rect 2955 16836 2959 16892
rect 2895 16832 2959 16836
rect 2975 16892 3039 16896
rect 2975 16836 2979 16892
rect 2979 16836 3035 16892
rect 3035 16836 3039 16892
rect 2975 16832 3039 16836
rect 3055 16892 3119 16896
rect 3055 16836 3059 16892
rect 3059 16836 3115 16892
rect 3115 16836 3119 16892
rect 3055 16832 3119 16836
rect 6541 16892 6605 16896
rect 6541 16836 6545 16892
rect 6545 16836 6601 16892
rect 6601 16836 6605 16892
rect 6541 16832 6605 16836
rect 6621 16892 6685 16896
rect 6621 16836 6625 16892
rect 6625 16836 6681 16892
rect 6681 16836 6685 16892
rect 6621 16832 6685 16836
rect 6701 16892 6765 16896
rect 6701 16836 6705 16892
rect 6705 16836 6761 16892
rect 6761 16836 6765 16892
rect 6701 16832 6765 16836
rect 6781 16892 6845 16896
rect 6781 16836 6785 16892
rect 6785 16836 6841 16892
rect 6841 16836 6845 16892
rect 6781 16832 6845 16836
rect 10267 16892 10331 16896
rect 10267 16836 10271 16892
rect 10271 16836 10327 16892
rect 10327 16836 10331 16892
rect 10267 16832 10331 16836
rect 10347 16892 10411 16896
rect 10347 16836 10351 16892
rect 10351 16836 10407 16892
rect 10407 16836 10411 16892
rect 10347 16832 10411 16836
rect 10427 16892 10491 16896
rect 10427 16836 10431 16892
rect 10431 16836 10487 16892
rect 10487 16836 10491 16892
rect 10427 16832 10491 16836
rect 10507 16892 10571 16896
rect 10507 16836 10511 16892
rect 10511 16836 10567 16892
rect 10567 16836 10571 16892
rect 10507 16832 10571 16836
rect 13993 16892 14057 16896
rect 13993 16836 13997 16892
rect 13997 16836 14053 16892
rect 14053 16836 14057 16892
rect 13993 16832 14057 16836
rect 14073 16892 14137 16896
rect 14073 16836 14077 16892
rect 14077 16836 14133 16892
rect 14133 16836 14137 16892
rect 14073 16832 14137 16836
rect 14153 16892 14217 16896
rect 14153 16836 14157 16892
rect 14157 16836 14213 16892
rect 14213 16836 14217 16892
rect 14153 16832 14217 16836
rect 14233 16892 14297 16896
rect 14233 16836 14237 16892
rect 14237 16836 14293 16892
rect 14293 16836 14297 16892
rect 14233 16832 14297 16836
rect 3475 16348 3539 16352
rect 3475 16292 3479 16348
rect 3479 16292 3535 16348
rect 3535 16292 3539 16348
rect 3475 16288 3539 16292
rect 3555 16348 3619 16352
rect 3555 16292 3559 16348
rect 3559 16292 3615 16348
rect 3615 16292 3619 16348
rect 3555 16288 3619 16292
rect 3635 16348 3699 16352
rect 3635 16292 3639 16348
rect 3639 16292 3695 16348
rect 3695 16292 3699 16348
rect 3635 16288 3699 16292
rect 3715 16348 3779 16352
rect 3715 16292 3719 16348
rect 3719 16292 3775 16348
rect 3775 16292 3779 16348
rect 3715 16288 3779 16292
rect 7201 16348 7265 16352
rect 7201 16292 7205 16348
rect 7205 16292 7261 16348
rect 7261 16292 7265 16348
rect 7201 16288 7265 16292
rect 7281 16348 7345 16352
rect 7281 16292 7285 16348
rect 7285 16292 7341 16348
rect 7341 16292 7345 16348
rect 7281 16288 7345 16292
rect 7361 16348 7425 16352
rect 7361 16292 7365 16348
rect 7365 16292 7421 16348
rect 7421 16292 7425 16348
rect 7361 16288 7425 16292
rect 7441 16348 7505 16352
rect 7441 16292 7445 16348
rect 7445 16292 7501 16348
rect 7501 16292 7505 16348
rect 7441 16288 7505 16292
rect 10927 16348 10991 16352
rect 10927 16292 10931 16348
rect 10931 16292 10987 16348
rect 10987 16292 10991 16348
rect 10927 16288 10991 16292
rect 11007 16348 11071 16352
rect 11007 16292 11011 16348
rect 11011 16292 11067 16348
rect 11067 16292 11071 16348
rect 11007 16288 11071 16292
rect 11087 16348 11151 16352
rect 11087 16292 11091 16348
rect 11091 16292 11147 16348
rect 11147 16292 11151 16348
rect 11087 16288 11151 16292
rect 11167 16348 11231 16352
rect 11167 16292 11171 16348
rect 11171 16292 11227 16348
rect 11227 16292 11231 16348
rect 11167 16288 11231 16292
rect 14653 16348 14717 16352
rect 14653 16292 14657 16348
rect 14657 16292 14713 16348
rect 14713 16292 14717 16348
rect 14653 16288 14717 16292
rect 14733 16348 14797 16352
rect 14733 16292 14737 16348
rect 14737 16292 14793 16348
rect 14793 16292 14797 16348
rect 14733 16288 14797 16292
rect 14813 16348 14877 16352
rect 14813 16292 14817 16348
rect 14817 16292 14873 16348
rect 14873 16292 14877 16348
rect 14813 16288 14877 16292
rect 14893 16348 14957 16352
rect 14893 16292 14897 16348
rect 14897 16292 14953 16348
rect 14953 16292 14957 16348
rect 14893 16288 14957 16292
rect 2815 15804 2879 15808
rect 2815 15748 2819 15804
rect 2819 15748 2875 15804
rect 2875 15748 2879 15804
rect 2815 15744 2879 15748
rect 2895 15804 2959 15808
rect 2895 15748 2899 15804
rect 2899 15748 2955 15804
rect 2955 15748 2959 15804
rect 2895 15744 2959 15748
rect 2975 15804 3039 15808
rect 2975 15748 2979 15804
rect 2979 15748 3035 15804
rect 3035 15748 3039 15804
rect 2975 15744 3039 15748
rect 3055 15804 3119 15808
rect 3055 15748 3059 15804
rect 3059 15748 3115 15804
rect 3115 15748 3119 15804
rect 3055 15744 3119 15748
rect 6541 15804 6605 15808
rect 6541 15748 6545 15804
rect 6545 15748 6601 15804
rect 6601 15748 6605 15804
rect 6541 15744 6605 15748
rect 6621 15804 6685 15808
rect 6621 15748 6625 15804
rect 6625 15748 6681 15804
rect 6681 15748 6685 15804
rect 6621 15744 6685 15748
rect 6701 15804 6765 15808
rect 6701 15748 6705 15804
rect 6705 15748 6761 15804
rect 6761 15748 6765 15804
rect 6701 15744 6765 15748
rect 6781 15804 6845 15808
rect 6781 15748 6785 15804
rect 6785 15748 6841 15804
rect 6841 15748 6845 15804
rect 6781 15744 6845 15748
rect 10267 15804 10331 15808
rect 10267 15748 10271 15804
rect 10271 15748 10327 15804
rect 10327 15748 10331 15804
rect 10267 15744 10331 15748
rect 10347 15804 10411 15808
rect 10347 15748 10351 15804
rect 10351 15748 10407 15804
rect 10407 15748 10411 15804
rect 10347 15744 10411 15748
rect 10427 15804 10491 15808
rect 10427 15748 10431 15804
rect 10431 15748 10487 15804
rect 10487 15748 10491 15804
rect 10427 15744 10491 15748
rect 10507 15804 10571 15808
rect 10507 15748 10511 15804
rect 10511 15748 10567 15804
rect 10567 15748 10571 15804
rect 10507 15744 10571 15748
rect 13993 15804 14057 15808
rect 13993 15748 13997 15804
rect 13997 15748 14053 15804
rect 14053 15748 14057 15804
rect 13993 15744 14057 15748
rect 14073 15804 14137 15808
rect 14073 15748 14077 15804
rect 14077 15748 14133 15804
rect 14133 15748 14137 15804
rect 14073 15744 14137 15748
rect 14153 15804 14217 15808
rect 14153 15748 14157 15804
rect 14157 15748 14213 15804
rect 14213 15748 14217 15804
rect 14153 15744 14217 15748
rect 14233 15804 14297 15808
rect 14233 15748 14237 15804
rect 14237 15748 14293 15804
rect 14293 15748 14297 15804
rect 14233 15744 14297 15748
rect 3475 15260 3539 15264
rect 3475 15204 3479 15260
rect 3479 15204 3535 15260
rect 3535 15204 3539 15260
rect 3475 15200 3539 15204
rect 3555 15260 3619 15264
rect 3555 15204 3559 15260
rect 3559 15204 3615 15260
rect 3615 15204 3619 15260
rect 3555 15200 3619 15204
rect 3635 15260 3699 15264
rect 3635 15204 3639 15260
rect 3639 15204 3695 15260
rect 3695 15204 3699 15260
rect 3635 15200 3699 15204
rect 3715 15260 3779 15264
rect 3715 15204 3719 15260
rect 3719 15204 3775 15260
rect 3775 15204 3779 15260
rect 3715 15200 3779 15204
rect 7201 15260 7265 15264
rect 7201 15204 7205 15260
rect 7205 15204 7261 15260
rect 7261 15204 7265 15260
rect 7201 15200 7265 15204
rect 7281 15260 7345 15264
rect 7281 15204 7285 15260
rect 7285 15204 7341 15260
rect 7341 15204 7345 15260
rect 7281 15200 7345 15204
rect 7361 15260 7425 15264
rect 7361 15204 7365 15260
rect 7365 15204 7421 15260
rect 7421 15204 7425 15260
rect 7361 15200 7425 15204
rect 7441 15260 7505 15264
rect 7441 15204 7445 15260
rect 7445 15204 7501 15260
rect 7501 15204 7505 15260
rect 7441 15200 7505 15204
rect 10927 15260 10991 15264
rect 10927 15204 10931 15260
rect 10931 15204 10987 15260
rect 10987 15204 10991 15260
rect 10927 15200 10991 15204
rect 11007 15260 11071 15264
rect 11007 15204 11011 15260
rect 11011 15204 11067 15260
rect 11067 15204 11071 15260
rect 11007 15200 11071 15204
rect 11087 15260 11151 15264
rect 11087 15204 11091 15260
rect 11091 15204 11147 15260
rect 11147 15204 11151 15260
rect 11087 15200 11151 15204
rect 11167 15260 11231 15264
rect 11167 15204 11171 15260
rect 11171 15204 11227 15260
rect 11227 15204 11231 15260
rect 11167 15200 11231 15204
rect 14653 15260 14717 15264
rect 14653 15204 14657 15260
rect 14657 15204 14713 15260
rect 14713 15204 14717 15260
rect 14653 15200 14717 15204
rect 14733 15260 14797 15264
rect 14733 15204 14737 15260
rect 14737 15204 14793 15260
rect 14793 15204 14797 15260
rect 14733 15200 14797 15204
rect 14813 15260 14877 15264
rect 14813 15204 14817 15260
rect 14817 15204 14873 15260
rect 14873 15204 14877 15260
rect 14813 15200 14877 15204
rect 14893 15260 14957 15264
rect 14893 15204 14897 15260
rect 14897 15204 14953 15260
rect 14953 15204 14957 15260
rect 14893 15200 14957 15204
rect 2815 14716 2879 14720
rect 2815 14660 2819 14716
rect 2819 14660 2875 14716
rect 2875 14660 2879 14716
rect 2815 14656 2879 14660
rect 2895 14716 2959 14720
rect 2895 14660 2899 14716
rect 2899 14660 2955 14716
rect 2955 14660 2959 14716
rect 2895 14656 2959 14660
rect 2975 14716 3039 14720
rect 2975 14660 2979 14716
rect 2979 14660 3035 14716
rect 3035 14660 3039 14716
rect 2975 14656 3039 14660
rect 3055 14716 3119 14720
rect 3055 14660 3059 14716
rect 3059 14660 3115 14716
rect 3115 14660 3119 14716
rect 3055 14656 3119 14660
rect 6541 14716 6605 14720
rect 6541 14660 6545 14716
rect 6545 14660 6601 14716
rect 6601 14660 6605 14716
rect 6541 14656 6605 14660
rect 6621 14716 6685 14720
rect 6621 14660 6625 14716
rect 6625 14660 6681 14716
rect 6681 14660 6685 14716
rect 6621 14656 6685 14660
rect 6701 14716 6765 14720
rect 6701 14660 6705 14716
rect 6705 14660 6761 14716
rect 6761 14660 6765 14716
rect 6701 14656 6765 14660
rect 6781 14716 6845 14720
rect 6781 14660 6785 14716
rect 6785 14660 6841 14716
rect 6841 14660 6845 14716
rect 6781 14656 6845 14660
rect 10267 14716 10331 14720
rect 10267 14660 10271 14716
rect 10271 14660 10327 14716
rect 10327 14660 10331 14716
rect 10267 14656 10331 14660
rect 10347 14716 10411 14720
rect 10347 14660 10351 14716
rect 10351 14660 10407 14716
rect 10407 14660 10411 14716
rect 10347 14656 10411 14660
rect 10427 14716 10491 14720
rect 10427 14660 10431 14716
rect 10431 14660 10487 14716
rect 10487 14660 10491 14716
rect 10427 14656 10491 14660
rect 10507 14716 10571 14720
rect 10507 14660 10511 14716
rect 10511 14660 10567 14716
rect 10567 14660 10571 14716
rect 10507 14656 10571 14660
rect 13993 14716 14057 14720
rect 13993 14660 13997 14716
rect 13997 14660 14053 14716
rect 14053 14660 14057 14716
rect 13993 14656 14057 14660
rect 14073 14716 14137 14720
rect 14073 14660 14077 14716
rect 14077 14660 14133 14716
rect 14133 14660 14137 14716
rect 14073 14656 14137 14660
rect 14153 14716 14217 14720
rect 14153 14660 14157 14716
rect 14157 14660 14213 14716
rect 14213 14660 14217 14716
rect 14153 14656 14217 14660
rect 14233 14716 14297 14720
rect 14233 14660 14237 14716
rect 14237 14660 14293 14716
rect 14293 14660 14297 14716
rect 14233 14656 14297 14660
rect 3475 14172 3539 14176
rect 3475 14116 3479 14172
rect 3479 14116 3535 14172
rect 3535 14116 3539 14172
rect 3475 14112 3539 14116
rect 3555 14172 3619 14176
rect 3555 14116 3559 14172
rect 3559 14116 3615 14172
rect 3615 14116 3619 14172
rect 3555 14112 3619 14116
rect 3635 14172 3699 14176
rect 3635 14116 3639 14172
rect 3639 14116 3695 14172
rect 3695 14116 3699 14172
rect 3635 14112 3699 14116
rect 3715 14172 3779 14176
rect 3715 14116 3719 14172
rect 3719 14116 3775 14172
rect 3775 14116 3779 14172
rect 3715 14112 3779 14116
rect 7201 14172 7265 14176
rect 7201 14116 7205 14172
rect 7205 14116 7261 14172
rect 7261 14116 7265 14172
rect 7201 14112 7265 14116
rect 7281 14172 7345 14176
rect 7281 14116 7285 14172
rect 7285 14116 7341 14172
rect 7341 14116 7345 14172
rect 7281 14112 7345 14116
rect 7361 14172 7425 14176
rect 7361 14116 7365 14172
rect 7365 14116 7421 14172
rect 7421 14116 7425 14172
rect 7361 14112 7425 14116
rect 7441 14172 7505 14176
rect 7441 14116 7445 14172
rect 7445 14116 7501 14172
rect 7501 14116 7505 14172
rect 7441 14112 7505 14116
rect 10927 14172 10991 14176
rect 10927 14116 10931 14172
rect 10931 14116 10987 14172
rect 10987 14116 10991 14172
rect 10927 14112 10991 14116
rect 11007 14172 11071 14176
rect 11007 14116 11011 14172
rect 11011 14116 11067 14172
rect 11067 14116 11071 14172
rect 11007 14112 11071 14116
rect 11087 14172 11151 14176
rect 11087 14116 11091 14172
rect 11091 14116 11147 14172
rect 11147 14116 11151 14172
rect 11087 14112 11151 14116
rect 11167 14172 11231 14176
rect 11167 14116 11171 14172
rect 11171 14116 11227 14172
rect 11227 14116 11231 14172
rect 11167 14112 11231 14116
rect 14653 14172 14717 14176
rect 14653 14116 14657 14172
rect 14657 14116 14713 14172
rect 14713 14116 14717 14172
rect 14653 14112 14717 14116
rect 14733 14172 14797 14176
rect 14733 14116 14737 14172
rect 14737 14116 14793 14172
rect 14793 14116 14797 14172
rect 14733 14112 14797 14116
rect 14813 14172 14877 14176
rect 14813 14116 14817 14172
rect 14817 14116 14873 14172
rect 14873 14116 14877 14172
rect 14813 14112 14877 14116
rect 14893 14172 14957 14176
rect 14893 14116 14897 14172
rect 14897 14116 14953 14172
rect 14953 14116 14957 14172
rect 14893 14112 14957 14116
rect 2815 13628 2879 13632
rect 2815 13572 2819 13628
rect 2819 13572 2875 13628
rect 2875 13572 2879 13628
rect 2815 13568 2879 13572
rect 2895 13628 2959 13632
rect 2895 13572 2899 13628
rect 2899 13572 2955 13628
rect 2955 13572 2959 13628
rect 2895 13568 2959 13572
rect 2975 13628 3039 13632
rect 2975 13572 2979 13628
rect 2979 13572 3035 13628
rect 3035 13572 3039 13628
rect 2975 13568 3039 13572
rect 3055 13628 3119 13632
rect 3055 13572 3059 13628
rect 3059 13572 3115 13628
rect 3115 13572 3119 13628
rect 3055 13568 3119 13572
rect 6541 13628 6605 13632
rect 6541 13572 6545 13628
rect 6545 13572 6601 13628
rect 6601 13572 6605 13628
rect 6541 13568 6605 13572
rect 6621 13628 6685 13632
rect 6621 13572 6625 13628
rect 6625 13572 6681 13628
rect 6681 13572 6685 13628
rect 6621 13568 6685 13572
rect 6701 13628 6765 13632
rect 6701 13572 6705 13628
rect 6705 13572 6761 13628
rect 6761 13572 6765 13628
rect 6701 13568 6765 13572
rect 6781 13628 6845 13632
rect 6781 13572 6785 13628
rect 6785 13572 6841 13628
rect 6841 13572 6845 13628
rect 6781 13568 6845 13572
rect 10267 13628 10331 13632
rect 10267 13572 10271 13628
rect 10271 13572 10327 13628
rect 10327 13572 10331 13628
rect 10267 13568 10331 13572
rect 10347 13628 10411 13632
rect 10347 13572 10351 13628
rect 10351 13572 10407 13628
rect 10407 13572 10411 13628
rect 10347 13568 10411 13572
rect 10427 13628 10491 13632
rect 10427 13572 10431 13628
rect 10431 13572 10487 13628
rect 10487 13572 10491 13628
rect 10427 13568 10491 13572
rect 10507 13628 10571 13632
rect 10507 13572 10511 13628
rect 10511 13572 10567 13628
rect 10567 13572 10571 13628
rect 10507 13568 10571 13572
rect 13993 13628 14057 13632
rect 13993 13572 13997 13628
rect 13997 13572 14053 13628
rect 14053 13572 14057 13628
rect 13993 13568 14057 13572
rect 14073 13628 14137 13632
rect 14073 13572 14077 13628
rect 14077 13572 14133 13628
rect 14133 13572 14137 13628
rect 14073 13568 14137 13572
rect 14153 13628 14217 13632
rect 14153 13572 14157 13628
rect 14157 13572 14213 13628
rect 14213 13572 14217 13628
rect 14153 13568 14217 13572
rect 14233 13628 14297 13632
rect 14233 13572 14237 13628
rect 14237 13572 14293 13628
rect 14293 13572 14297 13628
rect 14233 13568 14297 13572
rect 3475 13084 3539 13088
rect 3475 13028 3479 13084
rect 3479 13028 3535 13084
rect 3535 13028 3539 13084
rect 3475 13024 3539 13028
rect 3555 13084 3619 13088
rect 3555 13028 3559 13084
rect 3559 13028 3615 13084
rect 3615 13028 3619 13084
rect 3555 13024 3619 13028
rect 3635 13084 3699 13088
rect 3635 13028 3639 13084
rect 3639 13028 3695 13084
rect 3695 13028 3699 13084
rect 3635 13024 3699 13028
rect 3715 13084 3779 13088
rect 3715 13028 3719 13084
rect 3719 13028 3775 13084
rect 3775 13028 3779 13084
rect 3715 13024 3779 13028
rect 7201 13084 7265 13088
rect 7201 13028 7205 13084
rect 7205 13028 7261 13084
rect 7261 13028 7265 13084
rect 7201 13024 7265 13028
rect 7281 13084 7345 13088
rect 7281 13028 7285 13084
rect 7285 13028 7341 13084
rect 7341 13028 7345 13084
rect 7281 13024 7345 13028
rect 7361 13084 7425 13088
rect 7361 13028 7365 13084
rect 7365 13028 7421 13084
rect 7421 13028 7425 13084
rect 7361 13024 7425 13028
rect 7441 13084 7505 13088
rect 7441 13028 7445 13084
rect 7445 13028 7501 13084
rect 7501 13028 7505 13084
rect 7441 13024 7505 13028
rect 10927 13084 10991 13088
rect 10927 13028 10931 13084
rect 10931 13028 10987 13084
rect 10987 13028 10991 13084
rect 10927 13024 10991 13028
rect 11007 13084 11071 13088
rect 11007 13028 11011 13084
rect 11011 13028 11067 13084
rect 11067 13028 11071 13084
rect 11007 13024 11071 13028
rect 11087 13084 11151 13088
rect 11087 13028 11091 13084
rect 11091 13028 11147 13084
rect 11147 13028 11151 13084
rect 11087 13024 11151 13028
rect 11167 13084 11231 13088
rect 11167 13028 11171 13084
rect 11171 13028 11227 13084
rect 11227 13028 11231 13084
rect 11167 13024 11231 13028
rect 14653 13084 14717 13088
rect 14653 13028 14657 13084
rect 14657 13028 14713 13084
rect 14713 13028 14717 13084
rect 14653 13024 14717 13028
rect 14733 13084 14797 13088
rect 14733 13028 14737 13084
rect 14737 13028 14793 13084
rect 14793 13028 14797 13084
rect 14733 13024 14797 13028
rect 14813 13084 14877 13088
rect 14813 13028 14817 13084
rect 14817 13028 14873 13084
rect 14873 13028 14877 13084
rect 14813 13024 14877 13028
rect 14893 13084 14957 13088
rect 14893 13028 14897 13084
rect 14897 13028 14953 13084
rect 14953 13028 14957 13084
rect 14893 13024 14957 13028
rect 2815 12540 2879 12544
rect 2815 12484 2819 12540
rect 2819 12484 2875 12540
rect 2875 12484 2879 12540
rect 2815 12480 2879 12484
rect 2895 12540 2959 12544
rect 2895 12484 2899 12540
rect 2899 12484 2955 12540
rect 2955 12484 2959 12540
rect 2895 12480 2959 12484
rect 2975 12540 3039 12544
rect 2975 12484 2979 12540
rect 2979 12484 3035 12540
rect 3035 12484 3039 12540
rect 2975 12480 3039 12484
rect 3055 12540 3119 12544
rect 3055 12484 3059 12540
rect 3059 12484 3115 12540
rect 3115 12484 3119 12540
rect 3055 12480 3119 12484
rect 6541 12540 6605 12544
rect 6541 12484 6545 12540
rect 6545 12484 6601 12540
rect 6601 12484 6605 12540
rect 6541 12480 6605 12484
rect 6621 12540 6685 12544
rect 6621 12484 6625 12540
rect 6625 12484 6681 12540
rect 6681 12484 6685 12540
rect 6621 12480 6685 12484
rect 6701 12540 6765 12544
rect 6701 12484 6705 12540
rect 6705 12484 6761 12540
rect 6761 12484 6765 12540
rect 6701 12480 6765 12484
rect 6781 12540 6845 12544
rect 6781 12484 6785 12540
rect 6785 12484 6841 12540
rect 6841 12484 6845 12540
rect 6781 12480 6845 12484
rect 10267 12540 10331 12544
rect 10267 12484 10271 12540
rect 10271 12484 10327 12540
rect 10327 12484 10331 12540
rect 10267 12480 10331 12484
rect 10347 12540 10411 12544
rect 10347 12484 10351 12540
rect 10351 12484 10407 12540
rect 10407 12484 10411 12540
rect 10347 12480 10411 12484
rect 10427 12540 10491 12544
rect 10427 12484 10431 12540
rect 10431 12484 10487 12540
rect 10487 12484 10491 12540
rect 10427 12480 10491 12484
rect 10507 12540 10571 12544
rect 10507 12484 10511 12540
rect 10511 12484 10567 12540
rect 10567 12484 10571 12540
rect 10507 12480 10571 12484
rect 13993 12540 14057 12544
rect 13993 12484 13997 12540
rect 13997 12484 14053 12540
rect 14053 12484 14057 12540
rect 13993 12480 14057 12484
rect 14073 12540 14137 12544
rect 14073 12484 14077 12540
rect 14077 12484 14133 12540
rect 14133 12484 14137 12540
rect 14073 12480 14137 12484
rect 14153 12540 14217 12544
rect 14153 12484 14157 12540
rect 14157 12484 14213 12540
rect 14213 12484 14217 12540
rect 14153 12480 14217 12484
rect 14233 12540 14297 12544
rect 14233 12484 14237 12540
rect 14237 12484 14293 12540
rect 14293 12484 14297 12540
rect 14233 12480 14297 12484
rect 3475 11996 3539 12000
rect 3475 11940 3479 11996
rect 3479 11940 3535 11996
rect 3535 11940 3539 11996
rect 3475 11936 3539 11940
rect 3555 11996 3619 12000
rect 3555 11940 3559 11996
rect 3559 11940 3615 11996
rect 3615 11940 3619 11996
rect 3555 11936 3619 11940
rect 3635 11996 3699 12000
rect 3635 11940 3639 11996
rect 3639 11940 3695 11996
rect 3695 11940 3699 11996
rect 3635 11936 3699 11940
rect 3715 11996 3779 12000
rect 3715 11940 3719 11996
rect 3719 11940 3775 11996
rect 3775 11940 3779 11996
rect 3715 11936 3779 11940
rect 7201 11996 7265 12000
rect 7201 11940 7205 11996
rect 7205 11940 7261 11996
rect 7261 11940 7265 11996
rect 7201 11936 7265 11940
rect 7281 11996 7345 12000
rect 7281 11940 7285 11996
rect 7285 11940 7341 11996
rect 7341 11940 7345 11996
rect 7281 11936 7345 11940
rect 7361 11996 7425 12000
rect 7361 11940 7365 11996
rect 7365 11940 7421 11996
rect 7421 11940 7425 11996
rect 7361 11936 7425 11940
rect 7441 11996 7505 12000
rect 7441 11940 7445 11996
rect 7445 11940 7501 11996
rect 7501 11940 7505 11996
rect 7441 11936 7505 11940
rect 10927 11996 10991 12000
rect 10927 11940 10931 11996
rect 10931 11940 10987 11996
rect 10987 11940 10991 11996
rect 10927 11936 10991 11940
rect 11007 11996 11071 12000
rect 11007 11940 11011 11996
rect 11011 11940 11067 11996
rect 11067 11940 11071 11996
rect 11007 11936 11071 11940
rect 11087 11996 11151 12000
rect 11087 11940 11091 11996
rect 11091 11940 11147 11996
rect 11147 11940 11151 11996
rect 11087 11936 11151 11940
rect 11167 11996 11231 12000
rect 11167 11940 11171 11996
rect 11171 11940 11227 11996
rect 11227 11940 11231 11996
rect 11167 11936 11231 11940
rect 14653 11996 14717 12000
rect 14653 11940 14657 11996
rect 14657 11940 14713 11996
rect 14713 11940 14717 11996
rect 14653 11936 14717 11940
rect 14733 11996 14797 12000
rect 14733 11940 14737 11996
rect 14737 11940 14793 11996
rect 14793 11940 14797 11996
rect 14733 11936 14797 11940
rect 14813 11996 14877 12000
rect 14813 11940 14817 11996
rect 14817 11940 14873 11996
rect 14873 11940 14877 11996
rect 14813 11936 14877 11940
rect 14893 11996 14957 12000
rect 14893 11940 14897 11996
rect 14897 11940 14953 11996
rect 14953 11940 14957 11996
rect 14893 11936 14957 11940
rect 2815 11452 2879 11456
rect 2815 11396 2819 11452
rect 2819 11396 2875 11452
rect 2875 11396 2879 11452
rect 2815 11392 2879 11396
rect 2895 11452 2959 11456
rect 2895 11396 2899 11452
rect 2899 11396 2955 11452
rect 2955 11396 2959 11452
rect 2895 11392 2959 11396
rect 2975 11452 3039 11456
rect 2975 11396 2979 11452
rect 2979 11396 3035 11452
rect 3035 11396 3039 11452
rect 2975 11392 3039 11396
rect 3055 11452 3119 11456
rect 3055 11396 3059 11452
rect 3059 11396 3115 11452
rect 3115 11396 3119 11452
rect 3055 11392 3119 11396
rect 6541 11452 6605 11456
rect 6541 11396 6545 11452
rect 6545 11396 6601 11452
rect 6601 11396 6605 11452
rect 6541 11392 6605 11396
rect 6621 11452 6685 11456
rect 6621 11396 6625 11452
rect 6625 11396 6681 11452
rect 6681 11396 6685 11452
rect 6621 11392 6685 11396
rect 6701 11452 6765 11456
rect 6701 11396 6705 11452
rect 6705 11396 6761 11452
rect 6761 11396 6765 11452
rect 6701 11392 6765 11396
rect 6781 11452 6845 11456
rect 6781 11396 6785 11452
rect 6785 11396 6841 11452
rect 6841 11396 6845 11452
rect 6781 11392 6845 11396
rect 10267 11452 10331 11456
rect 10267 11396 10271 11452
rect 10271 11396 10327 11452
rect 10327 11396 10331 11452
rect 10267 11392 10331 11396
rect 10347 11452 10411 11456
rect 10347 11396 10351 11452
rect 10351 11396 10407 11452
rect 10407 11396 10411 11452
rect 10347 11392 10411 11396
rect 10427 11452 10491 11456
rect 10427 11396 10431 11452
rect 10431 11396 10487 11452
rect 10487 11396 10491 11452
rect 10427 11392 10491 11396
rect 10507 11452 10571 11456
rect 10507 11396 10511 11452
rect 10511 11396 10567 11452
rect 10567 11396 10571 11452
rect 10507 11392 10571 11396
rect 13993 11452 14057 11456
rect 13993 11396 13997 11452
rect 13997 11396 14053 11452
rect 14053 11396 14057 11452
rect 13993 11392 14057 11396
rect 14073 11452 14137 11456
rect 14073 11396 14077 11452
rect 14077 11396 14133 11452
rect 14133 11396 14137 11452
rect 14073 11392 14137 11396
rect 14153 11452 14217 11456
rect 14153 11396 14157 11452
rect 14157 11396 14213 11452
rect 14213 11396 14217 11452
rect 14153 11392 14217 11396
rect 14233 11452 14297 11456
rect 14233 11396 14237 11452
rect 14237 11396 14293 11452
rect 14293 11396 14297 11452
rect 14233 11392 14297 11396
rect 3475 10908 3539 10912
rect 3475 10852 3479 10908
rect 3479 10852 3535 10908
rect 3535 10852 3539 10908
rect 3475 10848 3539 10852
rect 3555 10908 3619 10912
rect 3555 10852 3559 10908
rect 3559 10852 3615 10908
rect 3615 10852 3619 10908
rect 3555 10848 3619 10852
rect 3635 10908 3699 10912
rect 3635 10852 3639 10908
rect 3639 10852 3695 10908
rect 3695 10852 3699 10908
rect 3635 10848 3699 10852
rect 3715 10908 3779 10912
rect 3715 10852 3719 10908
rect 3719 10852 3775 10908
rect 3775 10852 3779 10908
rect 3715 10848 3779 10852
rect 7201 10908 7265 10912
rect 7201 10852 7205 10908
rect 7205 10852 7261 10908
rect 7261 10852 7265 10908
rect 7201 10848 7265 10852
rect 7281 10908 7345 10912
rect 7281 10852 7285 10908
rect 7285 10852 7341 10908
rect 7341 10852 7345 10908
rect 7281 10848 7345 10852
rect 7361 10908 7425 10912
rect 7361 10852 7365 10908
rect 7365 10852 7421 10908
rect 7421 10852 7425 10908
rect 7361 10848 7425 10852
rect 7441 10908 7505 10912
rect 7441 10852 7445 10908
rect 7445 10852 7501 10908
rect 7501 10852 7505 10908
rect 7441 10848 7505 10852
rect 10927 10908 10991 10912
rect 10927 10852 10931 10908
rect 10931 10852 10987 10908
rect 10987 10852 10991 10908
rect 10927 10848 10991 10852
rect 11007 10908 11071 10912
rect 11007 10852 11011 10908
rect 11011 10852 11067 10908
rect 11067 10852 11071 10908
rect 11007 10848 11071 10852
rect 11087 10908 11151 10912
rect 11087 10852 11091 10908
rect 11091 10852 11147 10908
rect 11147 10852 11151 10908
rect 11087 10848 11151 10852
rect 11167 10908 11231 10912
rect 11167 10852 11171 10908
rect 11171 10852 11227 10908
rect 11227 10852 11231 10908
rect 11167 10848 11231 10852
rect 14653 10908 14717 10912
rect 14653 10852 14657 10908
rect 14657 10852 14713 10908
rect 14713 10852 14717 10908
rect 14653 10848 14717 10852
rect 14733 10908 14797 10912
rect 14733 10852 14737 10908
rect 14737 10852 14793 10908
rect 14793 10852 14797 10908
rect 14733 10848 14797 10852
rect 14813 10908 14877 10912
rect 14813 10852 14817 10908
rect 14817 10852 14873 10908
rect 14873 10852 14877 10908
rect 14813 10848 14877 10852
rect 14893 10908 14957 10912
rect 14893 10852 14897 10908
rect 14897 10852 14953 10908
rect 14953 10852 14957 10908
rect 14893 10848 14957 10852
rect 2815 10364 2879 10368
rect 2815 10308 2819 10364
rect 2819 10308 2875 10364
rect 2875 10308 2879 10364
rect 2815 10304 2879 10308
rect 2895 10364 2959 10368
rect 2895 10308 2899 10364
rect 2899 10308 2955 10364
rect 2955 10308 2959 10364
rect 2895 10304 2959 10308
rect 2975 10364 3039 10368
rect 2975 10308 2979 10364
rect 2979 10308 3035 10364
rect 3035 10308 3039 10364
rect 2975 10304 3039 10308
rect 3055 10364 3119 10368
rect 3055 10308 3059 10364
rect 3059 10308 3115 10364
rect 3115 10308 3119 10364
rect 3055 10304 3119 10308
rect 6541 10364 6605 10368
rect 6541 10308 6545 10364
rect 6545 10308 6601 10364
rect 6601 10308 6605 10364
rect 6541 10304 6605 10308
rect 6621 10364 6685 10368
rect 6621 10308 6625 10364
rect 6625 10308 6681 10364
rect 6681 10308 6685 10364
rect 6621 10304 6685 10308
rect 6701 10364 6765 10368
rect 6701 10308 6705 10364
rect 6705 10308 6761 10364
rect 6761 10308 6765 10364
rect 6701 10304 6765 10308
rect 6781 10364 6845 10368
rect 6781 10308 6785 10364
rect 6785 10308 6841 10364
rect 6841 10308 6845 10364
rect 6781 10304 6845 10308
rect 10267 10364 10331 10368
rect 10267 10308 10271 10364
rect 10271 10308 10327 10364
rect 10327 10308 10331 10364
rect 10267 10304 10331 10308
rect 10347 10364 10411 10368
rect 10347 10308 10351 10364
rect 10351 10308 10407 10364
rect 10407 10308 10411 10364
rect 10347 10304 10411 10308
rect 10427 10364 10491 10368
rect 10427 10308 10431 10364
rect 10431 10308 10487 10364
rect 10487 10308 10491 10364
rect 10427 10304 10491 10308
rect 10507 10364 10571 10368
rect 10507 10308 10511 10364
rect 10511 10308 10567 10364
rect 10567 10308 10571 10364
rect 10507 10304 10571 10308
rect 13993 10364 14057 10368
rect 13993 10308 13997 10364
rect 13997 10308 14053 10364
rect 14053 10308 14057 10364
rect 13993 10304 14057 10308
rect 14073 10364 14137 10368
rect 14073 10308 14077 10364
rect 14077 10308 14133 10364
rect 14133 10308 14137 10364
rect 14073 10304 14137 10308
rect 14153 10364 14217 10368
rect 14153 10308 14157 10364
rect 14157 10308 14213 10364
rect 14213 10308 14217 10364
rect 14153 10304 14217 10308
rect 14233 10364 14297 10368
rect 14233 10308 14237 10364
rect 14237 10308 14293 10364
rect 14293 10308 14297 10364
rect 14233 10304 14297 10308
rect 3475 9820 3539 9824
rect 3475 9764 3479 9820
rect 3479 9764 3535 9820
rect 3535 9764 3539 9820
rect 3475 9760 3539 9764
rect 3555 9820 3619 9824
rect 3555 9764 3559 9820
rect 3559 9764 3615 9820
rect 3615 9764 3619 9820
rect 3555 9760 3619 9764
rect 3635 9820 3699 9824
rect 3635 9764 3639 9820
rect 3639 9764 3695 9820
rect 3695 9764 3699 9820
rect 3635 9760 3699 9764
rect 3715 9820 3779 9824
rect 3715 9764 3719 9820
rect 3719 9764 3775 9820
rect 3775 9764 3779 9820
rect 3715 9760 3779 9764
rect 7201 9820 7265 9824
rect 7201 9764 7205 9820
rect 7205 9764 7261 9820
rect 7261 9764 7265 9820
rect 7201 9760 7265 9764
rect 7281 9820 7345 9824
rect 7281 9764 7285 9820
rect 7285 9764 7341 9820
rect 7341 9764 7345 9820
rect 7281 9760 7345 9764
rect 7361 9820 7425 9824
rect 7361 9764 7365 9820
rect 7365 9764 7421 9820
rect 7421 9764 7425 9820
rect 7361 9760 7425 9764
rect 7441 9820 7505 9824
rect 7441 9764 7445 9820
rect 7445 9764 7501 9820
rect 7501 9764 7505 9820
rect 7441 9760 7505 9764
rect 10927 9820 10991 9824
rect 10927 9764 10931 9820
rect 10931 9764 10987 9820
rect 10987 9764 10991 9820
rect 10927 9760 10991 9764
rect 11007 9820 11071 9824
rect 11007 9764 11011 9820
rect 11011 9764 11067 9820
rect 11067 9764 11071 9820
rect 11007 9760 11071 9764
rect 11087 9820 11151 9824
rect 11087 9764 11091 9820
rect 11091 9764 11147 9820
rect 11147 9764 11151 9820
rect 11087 9760 11151 9764
rect 11167 9820 11231 9824
rect 11167 9764 11171 9820
rect 11171 9764 11227 9820
rect 11227 9764 11231 9820
rect 11167 9760 11231 9764
rect 14653 9820 14717 9824
rect 14653 9764 14657 9820
rect 14657 9764 14713 9820
rect 14713 9764 14717 9820
rect 14653 9760 14717 9764
rect 14733 9820 14797 9824
rect 14733 9764 14737 9820
rect 14737 9764 14793 9820
rect 14793 9764 14797 9820
rect 14733 9760 14797 9764
rect 14813 9820 14877 9824
rect 14813 9764 14817 9820
rect 14817 9764 14873 9820
rect 14873 9764 14877 9820
rect 14813 9760 14877 9764
rect 14893 9820 14957 9824
rect 14893 9764 14897 9820
rect 14897 9764 14953 9820
rect 14953 9764 14957 9820
rect 14893 9760 14957 9764
rect 2815 9276 2879 9280
rect 2815 9220 2819 9276
rect 2819 9220 2875 9276
rect 2875 9220 2879 9276
rect 2815 9216 2879 9220
rect 2895 9276 2959 9280
rect 2895 9220 2899 9276
rect 2899 9220 2955 9276
rect 2955 9220 2959 9276
rect 2895 9216 2959 9220
rect 2975 9276 3039 9280
rect 2975 9220 2979 9276
rect 2979 9220 3035 9276
rect 3035 9220 3039 9276
rect 2975 9216 3039 9220
rect 3055 9276 3119 9280
rect 3055 9220 3059 9276
rect 3059 9220 3115 9276
rect 3115 9220 3119 9276
rect 3055 9216 3119 9220
rect 6541 9276 6605 9280
rect 6541 9220 6545 9276
rect 6545 9220 6601 9276
rect 6601 9220 6605 9276
rect 6541 9216 6605 9220
rect 6621 9276 6685 9280
rect 6621 9220 6625 9276
rect 6625 9220 6681 9276
rect 6681 9220 6685 9276
rect 6621 9216 6685 9220
rect 6701 9276 6765 9280
rect 6701 9220 6705 9276
rect 6705 9220 6761 9276
rect 6761 9220 6765 9276
rect 6701 9216 6765 9220
rect 6781 9276 6845 9280
rect 6781 9220 6785 9276
rect 6785 9220 6841 9276
rect 6841 9220 6845 9276
rect 6781 9216 6845 9220
rect 10267 9276 10331 9280
rect 10267 9220 10271 9276
rect 10271 9220 10327 9276
rect 10327 9220 10331 9276
rect 10267 9216 10331 9220
rect 10347 9276 10411 9280
rect 10347 9220 10351 9276
rect 10351 9220 10407 9276
rect 10407 9220 10411 9276
rect 10347 9216 10411 9220
rect 10427 9276 10491 9280
rect 10427 9220 10431 9276
rect 10431 9220 10487 9276
rect 10487 9220 10491 9276
rect 10427 9216 10491 9220
rect 10507 9276 10571 9280
rect 10507 9220 10511 9276
rect 10511 9220 10567 9276
rect 10567 9220 10571 9276
rect 10507 9216 10571 9220
rect 13993 9276 14057 9280
rect 13993 9220 13997 9276
rect 13997 9220 14053 9276
rect 14053 9220 14057 9276
rect 13993 9216 14057 9220
rect 14073 9276 14137 9280
rect 14073 9220 14077 9276
rect 14077 9220 14133 9276
rect 14133 9220 14137 9276
rect 14073 9216 14137 9220
rect 14153 9276 14217 9280
rect 14153 9220 14157 9276
rect 14157 9220 14213 9276
rect 14213 9220 14217 9276
rect 14153 9216 14217 9220
rect 14233 9276 14297 9280
rect 14233 9220 14237 9276
rect 14237 9220 14293 9276
rect 14293 9220 14297 9276
rect 14233 9216 14297 9220
rect 3475 8732 3539 8736
rect 3475 8676 3479 8732
rect 3479 8676 3535 8732
rect 3535 8676 3539 8732
rect 3475 8672 3539 8676
rect 3555 8732 3619 8736
rect 3555 8676 3559 8732
rect 3559 8676 3615 8732
rect 3615 8676 3619 8732
rect 3555 8672 3619 8676
rect 3635 8732 3699 8736
rect 3635 8676 3639 8732
rect 3639 8676 3695 8732
rect 3695 8676 3699 8732
rect 3635 8672 3699 8676
rect 3715 8732 3779 8736
rect 3715 8676 3719 8732
rect 3719 8676 3775 8732
rect 3775 8676 3779 8732
rect 3715 8672 3779 8676
rect 7201 8732 7265 8736
rect 7201 8676 7205 8732
rect 7205 8676 7261 8732
rect 7261 8676 7265 8732
rect 7201 8672 7265 8676
rect 7281 8732 7345 8736
rect 7281 8676 7285 8732
rect 7285 8676 7341 8732
rect 7341 8676 7345 8732
rect 7281 8672 7345 8676
rect 7361 8732 7425 8736
rect 7361 8676 7365 8732
rect 7365 8676 7421 8732
rect 7421 8676 7425 8732
rect 7361 8672 7425 8676
rect 7441 8732 7505 8736
rect 7441 8676 7445 8732
rect 7445 8676 7501 8732
rect 7501 8676 7505 8732
rect 7441 8672 7505 8676
rect 10927 8732 10991 8736
rect 10927 8676 10931 8732
rect 10931 8676 10987 8732
rect 10987 8676 10991 8732
rect 10927 8672 10991 8676
rect 11007 8732 11071 8736
rect 11007 8676 11011 8732
rect 11011 8676 11067 8732
rect 11067 8676 11071 8732
rect 11007 8672 11071 8676
rect 11087 8732 11151 8736
rect 11087 8676 11091 8732
rect 11091 8676 11147 8732
rect 11147 8676 11151 8732
rect 11087 8672 11151 8676
rect 11167 8732 11231 8736
rect 11167 8676 11171 8732
rect 11171 8676 11227 8732
rect 11227 8676 11231 8732
rect 11167 8672 11231 8676
rect 14653 8732 14717 8736
rect 14653 8676 14657 8732
rect 14657 8676 14713 8732
rect 14713 8676 14717 8732
rect 14653 8672 14717 8676
rect 14733 8732 14797 8736
rect 14733 8676 14737 8732
rect 14737 8676 14793 8732
rect 14793 8676 14797 8732
rect 14733 8672 14797 8676
rect 14813 8732 14877 8736
rect 14813 8676 14817 8732
rect 14817 8676 14873 8732
rect 14873 8676 14877 8732
rect 14813 8672 14877 8676
rect 14893 8732 14957 8736
rect 14893 8676 14897 8732
rect 14897 8676 14953 8732
rect 14953 8676 14957 8732
rect 14893 8672 14957 8676
rect 2815 8188 2879 8192
rect 2815 8132 2819 8188
rect 2819 8132 2875 8188
rect 2875 8132 2879 8188
rect 2815 8128 2879 8132
rect 2895 8188 2959 8192
rect 2895 8132 2899 8188
rect 2899 8132 2955 8188
rect 2955 8132 2959 8188
rect 2895 8128 2959 8132
rect 2975 8188 3039 8192
rect 2975 8132 2979 8188
rect 2979 8132 3035 8188
rect 3035 8132 3039 8188
rect 2975 8128 3039 8132
rect 3055 8188 3119 8192
rect 3055 8132 3059 8188
rect 3059 8132 3115 8188
rect 3115 8132 3119 8188
rect 3055 8128 3119 8132
rect 6541 8188 6605 8192
rect 6541 8132 6545 8188
rect 6545 8132 6601 8188
rect 6601 8132 6605 8188
rect 6541 8128 6605 8132
rect 6621 8188 6685 8192
rect 6621 8132 6625 8188
rect 6625 8132 6681 8188
rect 6681 8132 6685 8188
rect 6621 8128 6685 8132
rect 6701 8188 6765 8192
rect 6701 8132 6705 8188
rect 6705 8132 6761 8188
rect 6761 8132 6765 8188
rect 6701 8128 6765 8132
rect 6781 8188 6845 8192
rect 6781 8132 6785 8188
rect 6785 8132 6841 8188
rect 6841 8132 6845 8188
rect 6781 8128 6845 8132
rect 10267 8188 10331 8192
rect 10267 8132 10271 8188
rect 10271 8132 10327 8188
rect 10327 8132 10331 8188
rect 10267 8128 10331 8132
rect 10347 8188 10411 8192
rect 10347 8132 10351 8188
rect 10351 8132 10407 8188
rect 10407 8132 10411 8188
rect 10347 8128 10411 8132
rect 10427 8188 10491 8192
rect 10427 8132 10431 8188
rect 10431 8132 10487 8188
rect 10487 8132 10491 8188
rect 10427 8128 10491 8132
rect 10507 8188 10571 8192
rect 10507 8132 10511 8188
rect 10511 8132 10567 8188
rect 10567 8132 10571 8188
rect 10507 8128 10571 8132
rect 13993 8188 14057 8192
rect 13993 8132 13997 8188
rect 13997 8132 14053 8188
rect 14053 8132 14057 8188
rect 13993 8128 14057 8132
rect 14073 8188 14137 8192
rect 14073 8132 14077 8188
rect 14077 8132 14133 8188
rect 14133 8132 14137 8188
rect 14073 8128 14137 8132
rect 14153 8188 14217 8192
rect 14153 8132 14157 8188
rect 14157 8132 14213 8188
rect 14213 8132 14217 8188
rect 14153 8128 14217 8132
rect 14233 8188 14297 8192
rect 14233 8132 14237 8188
rect 14237 8132 14293 8188
rect 14293 8132 14297 8188
rect 14233 8128 14297 8132
rect 3475 7644 3539 7648
rect 3475 7588 3479 7644
rect 3479 7588 3535 7644
rect 3535 7588 3539 7644
rect 3475 7584 3539 7588
rect 3555 7644 3619 7648
rect 3555 7588 3559 7644
rect 3559 7588 3615 7644
rect 3615 7588 3619 7644
rect 3555 7584 3619 7588
rect 3635 7644 3699 7648
rect 3635 7588 3639 7644
rect 3639 7588 3695 7644
rect 3695 7588 3699 7644
rect 3635 7584 3699 7588
rect 3715 7644 3779 7648
rect 3715 7588 3719 7644
rect 3719 7588 3775 7644
rect 3775 7588 3779 7644
rect 3715 7584 3779 7588
rect 7201 7644 7265 7648
rect 7201 7588 7205 7644
rect 7205 7588 7261 7644
rect 7261 7588 7265 7644
rect 7201 7584 7265 7588
rect 7281 7644 7345 7648
rect 7281 7588 7285 7644
rect 7285 7588 7341 7644
rect 7341 7588 7345 7644
rect 7281 7584 7345 7588
rect 7361 7644 7425 7648
rect 7361 7588 7365 7644
rect 7365 7588 7421 7644
rect 7421 7588 7425 7644
rect 7361 7584 7425 7588
rect 7441 7644 7505 7648
rect 7441 7588 7445 7644
rect 7445 7588 7501 7644
rect 7501 7588 7505 7644
rect 7441 7584 7505 7588
rect 10927 7644 10991 7648
rect 10927 7588 10931 7644
rect 10931 7588 10987 7644
rect 10987 7588 10991 7644
rect 10927 7584 10991 7588
rect 11007 7644 11071 7648
rect 11007 7588 11011 7644
rect 11011 7588 11067 7644
rect 11067 7588 11071 7644
rect 11007 7584 11071 7588
rect 11087 7644 11151 7648
rect 11087 7588 11091 7644
rect 11091 7588 11147 7644
rect 11147 7588 11151 7644
rect 11087 7584 11151 7588
rect 11167 7644 11231 7648
rect 11167 7588 11171 7644
rect 11171 7588 11227 7644
rect 11227 7588 11231 7644
rect 11167 7584 11231 7588
rect 14653 7644 14717 7648
rect 14653 7588 14657 7644
rect 14657 7588 14713 7644
rect 14713 7588 14717 7644
rect 14653 7584 14717 7588
rect 14733 7644 14797 7648
rect 14733 7588 14737 7644
rect 14737 7588 14793 7644
rect 14793 7588 14797 7644
rect 14733 7584 14797 7588
rect 14813 7644 14877 7648
rect 14813 7588 14817 7644
rect 14817 7588 14873 7644
rect 14873 7588 14877 7644
rect 14813 7584 14877 7588
rect 14893 7644 14957 7648
rect 14893 7588 14897 7644
rect 14897 7588 14953 7644
rect 14953 7588 14957 7644
rect 14893 7584 14957 7588
rect 2815 7100 2879 7104
rect 2815 7044 2819 7100
rect 2819 7044 2875 7100
rect 2875 7044 2879 7100
rect 2815 7040 2879 7044
rect 2895 7100 2959 7104
rect 2895 7044 2899 7100
rect 2899 7044 2955 7100
rect 2955 7044 2959 7100
rect 2895 7040 2959 7044
rect 2975 7100 3039 7104
rect 2975 7044 2979 7100
rect 2979 7044 3035 7100
rect 3035 7044 3039 7100
rect 2975 7040 3039 7044
rect 3055 7100 3119 7104
rect 3055 7044 3059 7100
rect 3059 7044 3115 7100
rect 3115 7044 3119 7100
rect 3055 7040 3119 7044
rect 6541 7100 6605 7104
rect 6541 7044 6545 7100
rect 6545 7044 6601 7100
rect 6601 7044 6605 7100
rect 6541 7040 6605 7044
rect 6621 7100 6685 7104
rect 6621 7044 6625 7100
rect 6625 7044 6681 7100
rect 6681 7044 6685 7100
rect 6621 7040 6685 7044
rect 6701 7100 6765 7104
rect 6701 7044 6705 7100
rect 6705 7044 6761 7100
rect 6761 7044 6765 7100
rect 6701 7040 6765 7044
rect 6781 7100 6845 7104
rect 6781 7044 6785 7100
rect 6785 7044 6841 7100
rect 6841 7044 6845 7100
rect 6781 7040 6845 7044
rect 10267 7100 10331 7104
rect 10267 7044 10271 7100
rect 10271 7044 10327 7100
rect 10327 7044 10331 7100
rect 10267 7040 10331 7044
rect 10347 7100 10411 7104
rect 10347 7044 10351 7100
rect 10351 7044 10407 7100
rect 10407 7044 10411 7100
rect 10347 7040 10411 7044
rect 10427 7100 10491 7104
rect 10427 7044 10431 7100
rect 10431 7044 10487 7100
rect 10487 7044 10491 7100
rect 10427 7040 10491 7044
rect 10507 7100 10571 7104
rect 10507 7044 10511 7100
rect 10511 7044 10567 7100
rect 10567 7044 10571 7100
rect 10507 7040 10571 7044
rect 13993 7100 14057 7104
rect 13993 7044 13997 7100
rect 13997 7044 14053 7100
rect 14053 7044 14057 7100
rect 13993 7040 14057 7044
rect 14073 7100 14137 7104
rect 14073 7044 14077 7100
rect 14077 7044 14133 7100
rect 14133 7044 14137 7100
rect 14073 7040 14137 7044
rect 14153 7100 14217 7104
rect 14153 7044 14157 7100
rect 14157 7044 14213 7100
rect 14213 7044 14217 7100
rect 14153 7040 14217 7044
rect 14233 7100 14297 7104
rect 14233 7044 14237 7100
rect 14237 7044 14293 7100
rect 14293 7044 14297 7100
rect 14233 7040 14297 7044
rect 3475 6556 3539 6560
rect 3475 6500 3479 6556
rect 3479 6500 3535 6556
rect 3535 6500 3539 6556
rect 3475 6496 3539 6500
rect 3555 6556 3619 6560
rect 3555 6500 3559 6556
rect 3559 6500 3615 6556
rect 3615 6500 3619 6556
rect 3555 6496 3619 6500
rect 3635 6556 3699 6560
rect 3635 6500 3639 6556
rect 3639 6500 3695 6556
rect 3695 6500 3699 6556
rect 3635 6496 3699 6500
rect 3715 6556 3779 6560
rect 3715 6500 3719 6556
rect 3719 6500 3775 6556
rect 3775 6500 3779 6556
rect 3715 6496 3779 6500
rect 7201 6556 7265 6560
rect 7201 6500 7205 6556
rect 7205 6500 7261 6556
rect 7261 6500 7265 6556
rect 7201 6496 7265 6500
rect 7281 6556 7345 6560
rect 7281 6500 7285 6556
rect 7285 6500 7341 6556
rect 7341 6500 7345 6556
rect 7281 6496 7345 6500
rect 7361 6556 7425 6560
rect 7361 6500 7365 6556
rect 7365 6500 7421 6556
rect 7421 6500 7425 6556
rect 7361 6496 7425 6500
rect 7441 6556 7505 6560
rect 7441 6500 7445 6556
rect 7445 6500 7501 6556
rect 7501 6500 7505 6556
rect 7441 6496 7505 6500
rect 10927 6556 10991 6560
rect 10927 6500 10931 6556
rect 10931 6500 10987 6556
rect 10987 6500 10991 6556
rect 10927 6496 10991 6500
rect 11007 6556 11071 6560
rect 11007 6500 11011 6556
rect 11011 6500 11067 6556
rect 11067 6500 11071 6556
rect 11007 6496 11071 6500
rect 11087 6556 11151 6560
rect 11087 6500 11091 6556
rect 11091 6500 11147 6556
rect 11147 6500 11151 6556
rect 11087 6496 11151 6500
rect 11167 6556 11231 6560
rect 11167 6500 11171 6556
rect 11171 6500 11227 6556
rect 11227 6500 11231 6556
rect 11167 6496 11231 6500
rect 14653 6556 14717 6560
rect 14653 6500 14657 6556
rect 14657 6500 14713 6556
rect 14713 6500 14717 6556
rect 14653 6496 14717 6500
rect 14733 6556 14797 6560
rect 14733 6500 14737 6556
rect 14737 6500 14793 6556
rect 14793 6500 14797 6556
rect 14733 6496 14797 6500
rect 14813 6556 14877 6560
rect 14813 6500 14817 6556
rect 14817 6500 14873 6556
rect 14873 6500 14877 6556
rect 14813 6496 14877 6500
rect 14893 6556 14957 6560
rect 14893 6500 14897 6556
rect 14897 6500 14953 6556
rect 14953 6500 14957 6556
rect 14893 6496 14957 6500
rect 2815 6012 2879 6016
rect 2815 5956 2819 6012
rect 2819 5956 2875 6012
rect 2875 5956 2879 6012
rect 2815 5952 2879 5956
rect 2895 6012 2959 6016
rect 2895 5956 2899 6012
rect 2899 5956 2955 6012
rect 2955 5956 2959 6012
rect 2895 5952 2959 5956
rect 2975 6012 3039 6016
rect 2975 5956 2979 6012
rect 2979 5956 3035 6012
rect 3035 5956 3039 6012
rect 2975 5952 3039 5956
rect 3055 6012 3119 6016
rect 3055 5956 3059 6012
rect 3059 5956 3115 6012
rect 3115 5956 3119 6012
rect 3055 5952 3119 5956
rect 6541 6012 6605 6016
rect 6541 5956 6545 6012
rect 6545 5956 6601 6012
rect 6601 5956 6605 6012
rect 6541 5952 6605 5956
rect 6621 6012 6685 6016
rect 6621 5956 6625 6012
rect 6625 5956 6681 6012
rect 6681 5956 6685 6012
rect 6621 5952 6685 5956
rect 6701 6012 6765 6016
rect 6701 5956 6705 6012
rect 6705 5956 6761 6012
rect 6761 5956 6765 6012
rect 6701 5952 6765 5956
rect 6781 6012 6845 6016
rect 6781 5956 6785 6012
rect 6785 5956 6841 6012
rect 6841 5956 6845 6012
rect 6781 5952 6845 5956
rect 10267 6012 10331 6016
rect 10267 5956 10271 6012
rect 10271 5956 10327 6012
rect 10327 5956 10331 6012
rect 10267 5952 10331 5956
rect 10347 6012 10411 6016
rect 10347 5956 10351 6012
rect 10351 5956 10407 6012
rect 10407 5956 10411 6012
rect 10347 5952 10411 5956
rect 10427 6012 10491 6016
rect 10427 5956 10431 6012
rect 10431 5956 10487 6012
rect 10487 5956 10491 6012
rect 10427 5952 10491 5956
rect 10507 6012 10571 6016
rect 10507 5956 10511 6012
rect 10511 5956 10567 6012
rect 10567 5956 10571 6012
rect 10507 5952 10571 5956
rect 13993 6012 14057 6016
rect 13993 5956 13997 6012
rect 13997 5956 14053 6012
rect 14053 5956 14057 6012
rect 13993 5952 14057 5956
rect 14073 6012 14137 6016
rect 14073 5956 14077 6012
rect 14077 5956 14133 6012
rect 14133 5956 14137 6012
rect 14073 5952 14137 5956
rect 14153 6012 14217 6016
rect 14153 5956 14157 6012
rect 14157 5956 14213 6012
rect 14213 5956 14217 6012
rect 14153 5952 14217 5956
rect 14233 6012 14297 6016
rect 14233 5956 14237 6012
rect 14237 5956 14293 6012
rect 14293 5956 14297 6012
rect 14233 5952 14297 5956
rect 3475 5468 3539 5472
rect 3475 5412 3479 5468
rect 3479 5412 3535 5468
rect 3535 5412 3539 5468
rect 3475 5408 3539 5412
rect 3555 5468 3619 5472
rect 3555 5412 3559 5468
rect 3559 5412 3615 5468
rect 3615 5412 3619 5468
rect 3555 5408 3619 5412
rect 3635 5468 3699 5472
rect 3635 5412 3639 5468
rect 3639 5412 3695 5468
rect 3695 5412 3699 5468
rect 3635 5408 3699 5412
rect 3715 5468 3779 5472
rect 3715 5412 3719 5468
rect 3719 5412 3775 5468
rect 3775 5412 3779 5468
rect 3715 5408 3779 5412
rect 7201 5468 7265 5472
rect 7201 5412 7205 5468
rect 7205 5412 7261 5468
rect 7261 5412 7265 5468
rect 7201 5408 7265 5412
rect 7281 5468 7345 5472
rect 7281 5412 7285 5468
rect 7285 5412 7341 5468
rect 7341 5412 7345 5468
rect 7281 5408 7345 5412
rect 7361 5468 7425 5472
rect 7361 5412 7365 5468
rect 7365 5412 7421 5468
rect 7421 5412 7425 5468
rect 7361 5408 7425 5412
rect 7441 5468 7505 5472
rect 7441 5412 7445 5468
rect 7445 5412 7501 5468
rect 7501 5412 7505 5468
rect 7441 5408 7505 5412
rect 10927 5468 10991 5472
rect 10927 5412 10931 5468
rect 10931 5412 10987 5468
rect 10987 5412 10991 5468
rect 10927 5408 10991 5412
rect 11007 5468 11071 5472
rect 11007 5412 11011 5468
rect 11011 5412 11067 5468
rect 11067 5412 11071 5468
rect 11007 5408 11071 5412
rect 11087 5468 11151 5472
rect 11087 5412 11091 5468
rect 11091 5412 11147 5468
rect 11147 5412 11151 5468
rect 11087 5408 11151 5412
rect 11167 5468 11231 5472
rect 11167 5412 11171 5468
rect 11171 5412 11227 5468
rect 11227 5412 11231 5468
rect 11167 5408 11231 5412
rect 14653 5468 14717 5472
rect 14653 5412 14657 5468
rect 14657 5412 14713 5468
rect 14713 5412 14717 5468
rect 14653 5408 14717 5412
rect 14733 5468 14797 5472
rect 14733 5412 14737 5468
rect 14737 5412 14793 5468
rect 14793 5412 14797 5468
rect 14733 5408 14797 5412
rect 14813 5468 14877 5472
rect 14813 5412 14817 5468
rect 14817 5412 14873 5468
rect 14873 5412 14877 5468
rect 14813 5408 14877 5412
rect 14893 5468 14957 5472
rect 14893 5412 14897 5468
rect 14897 5412 14953 5468
rect 14953 5412 14957 5468
rect 14893 5408 14957 5412
rect 2815 4924 2879 4928
rect 2815 4868 2819 4924
rect 2819 4868 2875 4924
rect 2875 4868 2879 4924
rect 2815 4864 2879 4868
rect 2895 4924 2959 4928
rect 2895 4868 2899 4924
rect 2899 4868 2955 4924
rect 2955 4868 2959 4924
rect 2895 4864 2959 4868
rect 2975 4924 3039 4928
rect 2975 4868 2979 4924
rect 2979 4868 3035 4924
rect 3035 4868 3039 4924
rect 2975 4864 3039 4868
rect 3055 4924 3119 4928
rect 3055 4868 3059 4924
rect 3059 4868 3115 4924
rect 3115 4868 3119 4924
rect 3055 4864 3119 4868
rect 6541 4924 6605 4928
rect 6541 4868 6545 4924
rect 6545 4868 6601 4924
rect 6601 4868 6605 4924
rect 6541 4864 6605 4868
rect 6621 4924 6685 4928
rect 6621 4868 6625 4924
rect 6625 4868 6681 4924
rect 6681 4868 6685 4924
rect 6621 4864 6685 4868
rect 6701 4924 6765 4928
rect 6701 4868 6705 4924
rect 6705 4868 6761 4924
rect 6761 4868 6765 4924
rect 6701 4864 6765 4868
rect 6781 4924 6845 4928
rect 6781 4868 6785 4924
rect 6785 4868 6841 4924
rect 6841 4868 6845 4924
rect 6781 4864 6845 4868
rect 10267 4924 10331 4928
rect 10267 4868 10271 4924
rect 10271 4868 10327 4924
rect 10327 4868 10331 4924
rect 10267 4864 10331 4868
rect 10347 4924 10411 4928
rect 10347 4868 10351 4924
rect 10351 4868 10407 4924
rect 10407 4868 10411 4924
rect 10347 4864 10411 4868
rect 10427 4924 10491 4928
rect 10427 4868 10431 4924
rect 10431 4868 10487 4924
rect 10487 4868 10491 4924
rect 10427 4864 10491 4868
rect 10507 4924 10571 4928
rect 10507 4868 10511 4924
rect 10511 4868 10567 4924
rect 10567 4868 10571 4924
rect 10507 4864 10571 4868
rect 13993 4924 14057 4928
rect 13993 4868 13997 4924
rect 13997 4868 14053 4924
rect 14053 4868 14057 4924
rect 13993 4864 14057 4868
rect 14073 4924 14137 4928
rect 14073 4868 14077 4924
rect 14077 4868 14133 4924
rect 14133 4868 14137 4924
rect 14073 4864 14137 4868
rect 14153 4924 14217 4928
rect 14153 4868 14157 4924
rect 14157 4868 14213 4924
rect 14213 4868 14217 4924
rect 14153 4864 14217 4868
rect 14233 4924 14297 4928
rect 14233 4868 14237 4924
rect 14237 4868 14293 4924
rect 14293 4868 14297 4924
rect 14233 4864 14297 4868
rect 3475 4380 3539 4384
rect 3475 4324 3479 4380
rect 3479 4324 3535 4380
rect 3535 4324 3539 4380
rect 3475 4320 3539 4324
rect 3555 4380 3619 4384
rect 3555 4324 3559 4380
rect 3559 4324 3615 4380
rect 3615 4324 3619 4380
rect 3555 4320 3619 4324
rect 3635 4380 3699 4384
rect 3635 4324 3639 4380
rect 3639 4324 3695 4380
rect 3695 4324 3699 4380
rect 3635 4320 3699 4324
rect 3715 4380 3779 4384
rect 3715 4324 3719 4380
rect 3719 4324 3775 4380
rect 3775 4324 3779 4380
rect 3715 4320 3779 4324
rect 7201 4380 7265 4384
rect 7201 4324 7205 4380
rect 7205 4324 7261 4380
rect 7261 4324 7265 4380
rect 7201 4320 7265 4324
rect 7281 4380 7345 4384
rect 7281 4324 7285 4380
rect 7285 4324 7341 4380
rect 7341 4324 7345 4380
rect 7281 4320 7345 4324
rect 7361 4380 7425 4384
rect 7361 4324 7365 4380
rect 7365 4324 7421 4380
rect 7421 4324 7425 4380
rect 7361 4320 7425 4324
rect 7441 4380 7505 4384
rect 7441 4324 7445 4380
rect 7445 4324 7501 4380
rect 7501 4324 7505 4380
rect 7441 4320 7505 4324
rect 10927 4380 10991 4384
rect 10927 4324 10931 4380
rect 10931 4324 10987 4380
rect 10987 4324 10991 4380
rect 10927 4320 10991 4324
rect 11007 4380 11071 4384
rect 11007 4324 11011 4380
rect 11011 4324 11067 4380
rect 11067 4324 11071 4380
rect 11007 4320 11071 4324
rect 11087 4380 11151 4384
rect 11087 4324 11091 4380
rect 11091 4324 11147 4380
rect 11147 4324 11151 4380
rect 11087 4320 11151 4324
rect 11167 4380 11231 4384
rect 11167 4324 11171 4380
rect 11171 4324 11227 4380
rect 11227 4324 11231 4380
rect 11167 4320 11231 4324
rect 14653 4380 14717 4384
rect 14653 4324 14657 4380
rect 14657 4324 14713 4380
rect 14713 4324 14717 4380
rect 14653 4320 14717 4324
rect 14733 4380 14797 4384
rect 14733 4324 14737 4380
rect 14737 4324 14793 4380
rect 14793 4324 14797 4380
rect 14733 4320 14797 4324
rect 14813 4380 14877 4384
rect 14813 4324 14817 4380
rect 14817 4324 14873 4380
rect 14873 4324 14877 4380
rect 14813 4320 14877 4324
rect 14893 4380 14957 4384
rect 14893 4324 14897 4380
rect 14897 4324 14953 4380
rect 14953 4324 14957 4380
rect 14893 4320 14957 4324
rect 2815 3836 2879 3840
rect 2815 3780 2819 3836
rect 2819 3780 2875 3836
rect 2875 3780 2879 3836
rect 2815 3776 2879 3780
rect 2895 3836 2959 3840
rect 2895 3780 2899 3836
rect 2899 3780 2955 3836
rect 2955 3780 2959 3836
rect 2895 3776 2959 3780
rect 2975 3836 3039 3840
rect 2975 3780 2979 3836
rect 2979 3780 3035 3836
rect 3035 3780 3039 3836
rect 2975 3776 3039 3780
rect 3055 3836 3119 3840
rect 3055 3780 3059 3836
rect 3059 3780 3115 3836
rect 3115 3780 3119 3836
rect 3055 3776 3119 3780
rect 6541 3836 6605 3840
rect 6541 3780 6545 3836
rect 6545 3780 6601 3836
rect 6601 3780 6605 3836
rect 6541 3776 6605 3780
rect 6621 3836 6685 3840
rect 6621 3780 6625 3836
rect 6625 3780 6681 3836
rect 6681 3780 6685 3836
rect 6621 3776 6685 3780
rect 6701 3836 6765 3840
rect 6701 3780 6705 3836
rect 6705 3780 6761 3836
rect 6761 3780 6765 3836
rect 6701 3776 6765 3780
rect 6781 3836 6845 3840
rect 6781 3780 6785 3836
rect 6785 3780 6841 3836
rect 6841 3780 6845 3836
rect 6781 3776 6845 3780
rect 10267 3836 10331 3840
rect 10267 3780 10271 3836
rect 10271 3780 10327 3836
rect 10327 3780 10331 3836
rect 10267 3776 10331 3780
rect 10347 3836 10411 3840
rect 10347 3780 10351 3836
rect 10351 3780 10407 3836
rect 10407 3780 10411 3836
rect 10347 3776 10411 3780
rect 10427 3836 10491 3840
rect 10427 3780 10431 3836
rect 10431 3780 10487 3836
rect 10487 3780 10491 3836
rect 10427 3776 10491 3780
rect 10507 3836 10571 3840
rect 10507 3780 10511 3836
rect 10511 3780 10567 3836
rect 10567 3780 10571 3836
rect 10507 3776 10571 3780
rect 13993 3836 14057 3840
rect 13993 3780 13997 3836
rect 13997 3780 14053 3836
rect 14053 3780 14057 3836
rect 13993 3776 14057 3780
rect 14073 3836 14137 3840
rect 14073 3780 14077 3836
rect 14077 3780 14133 3836
rect 14133 3780 14137 3836
rect 14073 3776 14137 3780
rect 14153 3836 14217 3840
rect 14153 3780 14157 3836
rect 14157 3780 14213 3836
rect 14213 3780 14217 3836
rect 14153 3776 14217 3780
rect 14233 3836 14297 3840
rect 14233 3780 14237 3836
rect 14237 3780 14293 3836
rect 14293 3780 14297 3836
rect 14233 3776 14297 3780
rect 3475 3292 3539 3296
rect 3475 3236 3479 3292
rect 3479 3236 3535 3292
rect 3535 3236 3539 3292
rect 3475 3232 3539 3236
rect 3555 3292 3619 3296
rect 3555 3236 3559 3292
rect 3559 3236 3615 3292
rect 3615 3236 3619 3292
rect 3555 3232 3619 3236
rect 3635 3292 3699 3296
rect 3635 3236 3639 3292
rect 3639 3236 3695 3292
rect 3695 3236 3699 3292
rect 3635 3232 3699 3236
rect 3715 3292 3779 3296
rect 3715 3236 3719 3292
rect 3719 3236 3775 3292
rect 3775 3236 3779 3292
rect 3715 3232 3779 3236
rect 7201 3292 7265 3296
rect 7201 3236 7205 3292
rect 7205 3236 7261 3292
rect 7261 3236 7265 3292
rect 7201 3232 7265 3236
rect 7281 3292 7345 3296
rect 7281 3236 7285 3292
rect 7285 3236 7341 3292
rect 7341 3236 7345 3292
rect 7281 3232 7345 3236
rect 7361 3292 7425 3296
rect 7361 3236 7365 3292
rect 7365 3236 7421 3292
rect 7421 3236 7425 3292
rect 7361 3232 7425 3236
rect 7441 3292 7505 3296
rect 7441 3236 7445 3292
rect 7445 3236 7501 3292
rect 7501 3236 7505 3292
rect 7441 3232 7505 3236
rect 10927 3292 10991 3296
rect 10927 3236 10931 3292
rect 10931 3236 10987 3292
rect 10987 3236 10991 3292
rect 10927 3232 10991 3236
rect 11007 3292 11071 3296
rect 11007 3236 11011 3292
rect 11011 3236 11067 3292
rect 11067 3236 11071 3292
rect 11007 3232 11071 3236
rect 11087 3292 11151 3296
rect 11087 3236 11091 3292
rect 11091 3236 11147 3292
rect 11147 3236 11151 3292
rect 11087 3232 11151 3236
rect 11167 3292 11231 3296
rect 11167 3236 11171 3292
rect 11171 3236 11227 3292
rect 11227 3236 11231 3292
rect 11167 3232 11231 3236
rect 14653 3292 14717 3296
rect 14653 3236 14657 3292
rect 14657 3236 14713 3292
rect 14713 3236 14717 3292
rect 14653 3232 14717 3236
rect 14733 3292 14797 3296
rect 14733 3236 14737 3292
rect 14737 3236 14793 3292
rect 14793 3236 14797 3292
rect 14733 3232 14797 3236
rect 14813 3292 14877 3296
rect 14813 3236 14817 3292
rect 14817 3236 14873 3292
rect 14873 3236 14877 3292
rect 14813 3232 14877 3236
rect 14893 3292 14957 3296
rect 14893 3236 14897 3292
rect 14897 3236 14953 3292
rect 14953 3236 14957 3292
rect 14893 3232 14957 3236
rect 2815 2748 2879 2752
rect 2815 2692 2819 2748
rect 2819 2692 2875 2748
rect 2875 2692 2879 2748
rect 2815 2688 2879 2692
rect 2895 2748 2959 2752
rect 2895 2692 2899 2748
rect 2899 2692 2955 2748
rect 2955 2692 2959 2748
rect 2895 2688 2959 2692
rect 2975 2748 3039 2752
rect 2975 2692 2979 2748
rect 2979 2692 3035 2748
rect 3035 2692 3039 2748
rect 2975 2688 3039 2692
rect 3055 2748 3119 2752
rect 3055 2692 3059 2748
rect 3059 2692 3115 2748
rect 3115 2692 3119 2748
rect 3055 2688 3119 2692
rect 6541 2748 6605 2752
rect 6541 2692 6545 2748
rect 6545 2692 6601 2748
rect 6601 2692 6605 2748
rect 6541 2688 6605 2692
rect 6621 2748 6685 2752
rect 6621 2692 6625 2748
rect 6625 2692 6681 2748
rect 6681 2692 6685 2748
rect 6621 2688 6685 2692
rect 6701 2748 6765 2752
rect 6701 2692 6705 2748
rect 6705 2692 6761 2748
rect 6761 2692 6765 2748
rect 6701 2688 6765 2692
rect 6781 2748 6845 2752
rect 6781 2692 6785 2748
rect 6785 2692 6841 2748
rect 6841 2692 6845 2748
rect 6781 2688 6845 2692
rect 10267 2748 10331 2752
rect 10267 2692 10271 2748
rect 10271 2692 10327 2748
rect 10327 2692 10331 2748
rect 10267 2688 10331 2692
rect 10347 2748 10411 2752
rect 10347 2692 10351 2748
rect 10351 2692 10407 2748
rect 10407 2692 10411 2748
rect 10347 2688 10411 2692
rect 10427 2748 10491 2752
rect 10427 2692 10431 2748
rect 10431 2692 10487 2748
rect 10487 2692 10491 2748
rect 10427 2688 10491 2692
rect 10507 2748 10571 2752
rect 10507 2692 10511 2748
rect 10511 2692 10567 2748
rect 10567 2692 10571 2748
rect 10507 2688 10571 2692
rect 13993 2748 14057 2752
rect 13993 2692 13997 2748
rect 13997 2692 14053 2748
rect 14053 2692 14057 2748
rect 13993 2688 14057 2692
rect 14073 2748 14137 2752
rect 14073 2692 14077 2748
rect 14077 2692 14133 2748
rect 14133 2692 14137 2748
rect 14073 2688 14137 2692
rect 14153 2748 14217 2752
rect 14153 2692 14157 2748
rect 14157 2692 14213 2748
rect 14213 2692 14217 2748
rect 14153 2688 14217 2692
rect 14233 2748 14297 2752
rect 14233 2692 14237 2748
rect 14237 2692 14293 2748
rect 14293 2692 14297 2748
rect 14233 2688 14297 2692
rect 3475 2204 3539 2208
rect 3475 2148 3479 2204
rect 3479 2148 3535 2204
rect 3535 2148 3539 2204
rect 3475 2144 3539 2148
rect 3555 2204 3619 2208
rect 3555 2148 3559 2204
rect 3559 2148 3615 2204
rect 3615 2148 3619 2204
rect 3555 2144 3619 2148
rect 3635 2204 3699 2208
rect 3635 2148 3639 2204
rect 3639 2148 3695 2204
rect 3695 2148 3699 2204
rect 3635 2144 3699 2148
rect 3715 2204 3779 2208
rect 3715 2148 3719 2204
rect 3719 2148 3775 2204
rect 3775 2148 3779 2204
rect 3715 2144 3779 2148
rect 7201 2204 7265 2208
rect 7201 2148 7205 2204
rect 7205 2148 7261 2204
rect 7261 2148 7265 2204
rect 7201 2144 7265 2148
rect 7281 2204 7345 2208
rect 7281 2148 7285 2204
rect 7285 2148 7341 2204
rect 7341 2148 7345 2204
rect 7281 2144 7345 2148
rect 7361 2204 7425 2208
rect 7361 2148 7365 2204
rect 7365 2148 7421 2204
rect 7421 2148 7425 2204
rect 7361 2144 7425 2148
rect 7441 2204 7505 2208
rect 7441 2148 7445 2204
rect 7445 2148 7501 2204
rect 7501 2148 7505 2204
rect 7441 2144 7505 2148
rect 10927 2204 10991 2208
rect 10927 2148 10931 2204
rect 10931 2148 10987 2204
rect 10987 2148 10991 2204
rect 10927 2144 10991 2148
rect 11007 2204 11071 2208
rect 11007 2148 11011 2204
rect 11011 2148 11067 2204
rect 11067 2148 11071 2204
rect 11007 2144 11071 2148
rect 11087 2204 11151 2208
rect 11087 2148 11091 2204
rect 11091 2148 11147 2204
rect 11147 2148 11151 2204
rect 11087 2144 11151 2148
rect 11167 2204 11231 2208
rect 11167 2148 11171 2204
rect 11171 2148 11227 2204
rect 11227 2148 11231 2204
rect 11167 2144 11231 2148
rect 14653 2204 14717 2208
rect 14653 2148 14657 2204
rect 14657 2148 14713 2204
rect 14713 2148 14717 2204
rect 14653 2144 14717 2148
rect 14733 2204 14797 2208
rect 14733 2148 14737 2204
rect 14737 2148 14793 2204
rect 14793 2148 14797 2204
rect 14733 2144 14797 2148
rect 14813 2204 14877 2208
rect 14813 2148 14817 2204
rect 14817 2148 14873 2204
rect 14873 2148 14877 2204
rect 14813 2144 14877 2148
rect 14893 2204 14957 2208
rect 14893 2148 14897 2204
rect 14897 2148 14953 2204
rect 14953 2148 14957 2204
rect 14893 2144 14957 2148
<< metal4 >>
rect 2807 16896 3127 16912
rect 2807 16832 2815 16896
rect 2879 16832 2895 16896
rect 2959 16832 2975 16896
rect 3039 16832 3055 16896
rect 3119 16832 3127 16896
rect 2807 15808 3127 16832
rect 2807 15744 2815 15808
rect 2879 15744 2895 15808
rect 2959 15744 2975 15808
rect 3039 15744 3055 15808
rect 3119 15744 3127 15808
rect 2807 15146 3127 15744
rect 2807 14910 2849 15146
rect 3085 14910 3127 15146
rect 2807 14720 3127 14910
rect 2807 14656 2815 14720
rect 2879 14656 2895 14720
rect 2959 14656 2975 14720
rect 3039 14656 3055 14720
rect 3119 14656 3127 14720
rect 2807 13632 3127 14656
rect 2807 13568 2815 13632
rect 2879 13568 2895 13632
rect 2959 13568 2975 13632
rect 3039 13568 3055 13632
rect 3119 13568 3127 13632
rect 2807 12544 3127 13568
rect 2807 12480 2815 12544
rect 2879 12480 2895 12544
rect 2959 12480 2975 12544
rect 3039 12480 3055 12544
rect 3119 12480 3127 12544
rect 2807 11474 3127 12480
rect 2807 11456 2849 11474
rect 3085 11456 3127 11474
rect 2807 11392 2815 11456
rect 3119 11392 3127 11456
rect 2807 11238 2849 11392
rect 3085 11238 3127 11392
rect 2807 10368 3127 11238
rect 2807 10304 2815 10368
rect 2879 10304 2895 10368
rect 2959 10304 2975 10368
rect 3039 10304 3055 10368
rect 3119 10304 3127 10368
rect 2807 9280 3127 10304
rect 2807 9216 2815 9280
rect 2879 9216 2895 9280
rect 2959 9216 2975 9280
rect 3039 9216 3055 9280
rect 3119 9216 3127 9280
rect 2807 8192 3127 9216
rect 2807 8128 2815 8192
rect 2879 8128 2895 8192
rect 2959 8128 2975 8192
rect 3039 8128 3055 8192
rect 3119 8128 3127 8192
rect 2807 7802 3127 8128
rect 2807 7566 2849 7802
rect 3085 7566 3127 7802
rect 2807 7104 3127 7566
rect 2807 7040 2815 7104
rect 2879 7040 2895 7104
rect 2959 7040 2975 7104
rect 3039 7040 3055 7104
rect 3119 7040 3127 7104
rect 2807 6016 3127 7040
rect 2807 5952 2815 6016
rect 2879 5952 2895 6016
rect 2959 5952 2975 6016
rect 3039 5952 3055 6016
rect 3119 5952 3127 6016
rect 2807 4928 3127 5952
rect 2807 4864 2815 4928
rect 2879 4864 2895 4928
rect 2959 4864 2975 4928
rect 3039 4864 3055 4928
rect 3119 4864 3127 4928
rect 2807 4130 3127 4864
rect 2807 3894 2849 4130
rect 3085 3894 3127 4130
rect 2807 3840 3127 3894
rect 2807 3776 2815 3840
rect 2879 3776 2895 3840
rect 2959 3776 2975 3840
rect 3039 3776 3055 3840
rect 3119 3776 3127 3840
rect 2807 2752 3127 3776
rect 2807 2688 2815 2752
rect 2879 2688 2895 2752
rect 2959 2688 2975 2752
rect 3039 2688 3055 2752
rect 3119 2688 3127 2752
rect 2807 2128 3127 2688
rect 3467 16352 3787 16912
rect 3467 16288 3475 16352
rect 3539 16288 3555 16352
rect 3619 16288 3635 16352
rect 3699 16288 3715 16352
rect 3779 16288 3787 16352
rect 3467 15806 3787 16288
rect 3467 15570 3509 15806
rect 3745 15570 3787 15806
rect 3467 15264 3787 15570
rect 3467 15200 3475 15264
rect 3539 15200 3555 15264
rect 3619 15200 3635 15264
rect 3699 15200 3715 15264
rect 3779 15200 3787 15264
rect 3467 14176 3787 15200
rect 3467 14112 3475 14176
rect 3539 14112 3555 14176
rect 3619 14112 3635 14176
rect 3699 14112 3715 14176
rect 3779 14112 3787 14176
rect 3467 13088 3787 14112
rect 3467 13024 3475 13088
rect 3539 13024 3555 13088
rect 3619 13024 3635 13088
rect 3699 13024 3715 13088
rect 3779 13024 3787 13088
rect 3467 12134 3787 13024
rect 3467 12000 3509 12134
rect 3745 12000 3787 12134
rect 3467 11936 3475 12000
rect 3779 11936 3787 12000
rect 3467 11898 3509 11936
rect 3745 11898 3787 11936
rect 3467 10912 3787 11898
rect 3467 10848 3475 10912
rect 3539 10848 3555 10912
rect 3619 10848 3635 10912
rect 3699 10848 3715 10912
rect 3779 10848 3787 10912
rect 3467 9824 3787 10848
rect 3467 9760 3475 9824
rect 3539 9760 3555 9824
rect 3619 9760 3635 9824
rect 3699 9760 3715 9824
rect 3779 9760 3787 9824
rect 3467 8736 3787 9760
rect 3467 8672 3475 8736
rect 3539 8672 3555 8736
rect 3619 8672 3635 8736
rect 3699 8672 3715 8736
rect 3779 8672 3787 8736
rect 3467 8462 3787 8672
rect 3467 8226 3509 8462
rect 3745 8226 3787 8462
rect 3467 7648 3787 8226
rect 3467 7584 3475 7648
rect 3539 7584 3555 7648
rect 3619 7584 3635 7648
rect 3699 7584 3715 7648
rect 3779 7584 3787 7648
rect 3467 6560 3787 7584
rect 3467 6496 3475 6560
rect 3539 6496 3555 6560
rect 3619 6496 3635 6560
rect 3699 6496 3715 6560
rect 3779 6496 3787 6560
rect 3467 5472 3787 6496
rect 3467 5408 3475 5472
rect 3539 5408 3555 5472
rect 3619 5408 3635 5472
rect 3699 5408 3715 5472
rect 3779 5408 3787 5472
rect 3467 4790 3787 5408
rect 3467 4554 3509 4790
rect 3745 4554 3787 4790
rect 3467 4384 3787 4554
rect 3467 4320 3475 4384
rect 3539 4320 3555 4384
rect 3619 4320 3635 4384
rect 3699 4320 3715 4384
rect 3779 4320 3787 4384
rect 3467 3296 3787 4320
rect 3467 3232 3475 3296
rect 3539 3232 3555 3296
rect 3619 3232 3635 3296
rect 3699 3232 3715 3296
rect 3779 3232 3787 3296
rect 3467 2208 3787 3232
rect 3467 2144 3475 2208
rect 3539 2144 3555 2208
rect 3619 2144 3635 2208
rect 3699 2144 3715 2208
rect 3779 2144 3787 2208
rect 3467 2128 3787 2144
rect 6533 16896 6853 16912
rect 6533 16832 6541 16896
rect 6605 16832 6621 16896
rect 6685 16832 6701 16896
rect 6765 16832 6781 16896
rect 6845 16832 6853 16896
rect 6533 15808 6853 16832
rect 6533 15744 6541 15808
rect 6605 15744 6621 15808
rect 6685 15744 6701 15808
rect 6765 15744 6781 15808
rect 6845 15744 6853 15808
rect 6533 15146 6853 15744
rect 6533 14910 6575 15146
rect 6811 14910 6853 15146
rect 6533 14720 6853 14910
rect 6533 14656 6541 14720
rect 6605 14656 6621 14720
rect 6685 14656 6701 14720
rect 6765 14656 6781 14720
rect 6845 14656 6853 14720
rect 6533 13632 6853 14656
rect 6533 13568 6541 13632
rect 6605 13568 6621 13632
rect 6685 13568 6701 13632
rect 6765 13568 6781 13632
rect 6845 13568 6853 13632
rect 6533 12544 6853 13568
rect 6533 12480 6541 12544
rect 6605 12480 6621 12544
rect 6685 12480 6701 12544
rect 6765 12480 6781 12544
rect 6845 12480 6853 12544
rect 6533 11474 6853 12480
rect 6533 11456 6575 11474
rect 6811 11456 6853 11474
rect 6533 11392 6541 11456
rect 6845 11392 6853 11456
rect 6533 11238 6575 11392
rect 6811 11238 6853 11392
rect 6533 10368 6853 11238
rect 6533 10304 6541 10368
rect 6605 10304 6621 10368
rect 6685 10304 6701 10368
rect 6765 10304 6781 10368
rect 6845 10304 6853 10368
rect 6533 9280 6853 10304
rect 6533 9216 6541 9280
rect 6605 9216 6621 9280
rect 6685 9216 6701 9280
rect 6765 9216 6781 9280
rect 6845 9216 6853 9280
rect 6533 8192 6853 9216
rect 6533 8128 6541 8192
rect 6605 8128 6621 8192
rect 6685 8128 6701 8192
rect 6765 8128 6781 8192
rect 6845 8128 6853 8192
rect 6533 7802 6853 8128
rect 6533 7566 6575 7802
rect 6811 7566 6853 7802
rect 6533 7104 6853 7566
rect 6533 7040 6541 7104
rect 6605 7040 6621 7104
rect 6685 7040 6701 7104
rect 6765 7040 6781 7104
rect 6845 7040 6853 7104
rect 6533 6016 6853 7040
rect 6533 5952 6541 6016
rect 6605 5952 6621 6016
rect 6685 5952 6701 6016
rect 6765 5952 6781 6016
rect 6845 5952 6853 6016
rect 6533 4928 6853 5952
rect 6533 4864 6541 4928
rect 6605 4864 6621 4928
rect 6685 4864 6701 4928
rect 6765 4864 6781 4928
rect 6845 4864 6853 4928
rect 6533 4130 6853 4864
rect 6533 3894 6575 4130
rect 6811 3894 6853 4130
rect 6533 3840 6853 3894
rect 6533 3776 6541 3840
rect 6605 3776 6621 3840
rect 6685 3776 6701 3840
rect 6765 3776 6781 3840
rect 6845 3776 6853 3840
rect 6533 2752 6853 3776
rect 6533 2688 6541 2752
rect 6605 2688 6621 2752
rect 6685 2688 6701 2752
rect 6765 2688 6781 2752
rect 6845 2688 6853 2752
rect 6533 2128 6853 2688
rect 7193 16352 7513 16912
rect 7193 16288 7201 16352
rect 7265 16288 7281 16352
rect 7345 16288 7361 16352
rect 7425 16288 7441 16352
rect 7505 16288 7513 16352
rect 7193 15806 7513 16288
rect 7193 15570 7235 15806
rect 7471 15570 7513 15806
rect 7193 15264 7513 15570
rect 7193 15200 7201 15264
rect 7265 15200 7281 15264
rect 7345 15200 7361 15264
rect 7425 15200 7441 15264
rect 7505 15200 7513 15264
rect 7193 14176 7513 15200
rect 7193 14112 7201 14176
rect 7265 14112 7281 14176
rect 7345 14112 7361 14176
rect 7425 14112 7441 14176
rect 7505 14112 7513 14176
rect 7193 13088 7513 14112
rect 7193 13024 7201 13088
rect 7265 13024 7281 13088
rect 7345 13024 7361 13088
rect 7425 13024 7441 13088
rect 7505 13024 7513 13088
rect 7193 12134 7513 13024
rect 7193 12000 7235 12134
rect 7471 12000 7513 12134
rect 7193 11936 7201 12000
rect 7505 11936 7513 12000
rect 7193 11898 7235 11936
rect 7471 11898 7513 11936
rect 7193 10912 7513 11898
rect 7193 10848 7201 10912
rect 7265 10848 7281 10912
rect 7345 10848 7361 10912
rect 7425 10848 7441 10912
rect 7505 10848 7513 10912
rect 7193 9824 7513 10848
rect 7193 9760 7201 9824
rect 7265 9760 7281 9824
rect 7345 9760 7361 9824
rect 7425 9760 7441 9824
rect 7505 9760 7513 9824
rect 7193 8736 7513 9760
rect 7193 8672 7201 8736
rect 7265 8672 7281 8736
rect 7345 8672 7361 8736
rect 7425 8672 7441 8736
rect 7505 8672 7513 8736
rect 7193 8462 7513 8672
rect 7193 8226 7235 8462
rect 7471 8226 7513 8462
rect 7193 7648 7513 8226
rect 7193 7584 7201 7648
rect 7265 7584 7281 7648
rect 7345 7584 7361 7648
rect 7425 7584 7441 7648
rect 7505 7584 7513 7648
rect 7193 6560 7513 7584
rect 7193 6496 7201 6560
rect 7265 6496 7281 6560
rect 7345 6496 7361 6560
rect 7425 6496 7441 6560
rect 7505 6496 7513 6560
rect 7193 5472 7513 6496
rect 7193 5408 7201 5472
rect 7265 5408 7281 5472
rect 7345 5408 7361 5472
rect 7425 5408 7441 5472
rect 7505 5408 7513 5472
rect 7193 4790 7513 5408
rect 7193 4554 7235 4790
rect 7471 4554 7513 4790
rect 7193 4384 7513 4554
rect 7193 4320 7201 4384
rect 7265 4320 7281 4384
rect 7345 4320 7361 4384
rect 7425 4320 7441 4384
rect 7505 4320 7513 4384
rect 7193 3296 7513 4320
rect 7193 3232 7201 3296
rect 7265 3232 7281 3296
rect 7345 3232 7361 3296
rect 7425 3232 7441 3296
rect 7505 3232 7513 3296
rect 7193 2208 7513 3232
rect 7193 2144 7201 2208
rect 7265 2144 7281 2208
rect 7345 2144 7361 2208
rect 7425 2144 7441 2208
rect 7505 2144 7513 2208
rect 7193 2128 7513 2144
rect 10259 16896 10579 16912
rect 10259 16832 10267 16896
rect 10331 16832 10347 16896
rect 10411 16832 10427 16896
rect 10491 16832 10507 16896
rect 10571 16832 10579 16896
rect 10259 15808 10579 16832
rect 10259 15744 10267 15808
rect 10331 15744 10347 15808
rect 10411 15744 10427 15808
rect 10491 15744 10507 15808
rect 10571 15744 10579 15808
rect 10259 15146 10579 15744
rect 10259 14910 10301 15146
rect 10537 14910 10579 15146
rect 10259 14720 10579 14910
rect 10259 14656 10267 14720
rect 10331 14656 10347 14720
rect 10411 14656 10427 14720
rect 10491 14656 10507 14720
rect 10571 14656 10579 14720
rect 10259 13632 10579 14656
rect 10259 13568 10267 13632
rect 10331 13568 10347 13632
rect 10411 13568 10427 13632
rect 10491 13568 10507 13632
rect 10571 13568 10579 13632
rect 10259 12544 10579 13568
rect 10259 12480 10267 12544
rect 10331 12480 10347 12544
rect 10411 12480 10427 12544
rect 10491 12480 10507 12544
rect 10571 12480 10579 12544
rect 10259 11474 10579 12480
rect 10259 11456 10301 11474
rect 10537 11456 10579 11474
rect 10259 11392 10267 11456
rect 10571 11392 10579 11456
rect 10259 11238 10301 11392
rect 10537 11238 10579 11392
rect 10259 10368 10579 11238
rect 10259 10304 10267 10368
rect 10331 10304 10347 10368
rect 10411 10304 10427 10368
rect 10491 10304 10507 10368
rect 10571 10304 10579 10368
rect 10259 9280 10579 10304
rect 10259 9216 10267 9280
rect 10331 9216 10347 9280
rect 10411 9216 10427 9280
rect 10491 9216 10507 9280
rect 10571 9216 10579 9280
rect 10259 8192 10579 9216
rect 10259 8128 10267 8192
rect 10331 8128 10347 8192
rect 10411 8128 10427 8192
rect 10491 8128 10507 8192
rect 10571 8128 10579 8192
rect 10259 7802 10579 8128
rect 10259 7566 10301 7802
rect 10537 7566 10579 7802
rect 10259 7104 10579 7566
rect 10259 7040 10267 7104
rect 10331 7040 10347 7104
rect 10411 7040 10427 7104
rect 10491 7040 10507 7104
rect 10571 7040 10579 7104
rect 10259 6016 10579 7040
rect 10259 5952 10267 6016
rect 10331 5952 10347 6016
rect 10411 5952 10427 6016
rect 10491 5952 10507 6016
rect 10571 5952 10579 6016
rect 10259 4928 10579 5952
rect 10259 4864 10267 4928
rect 10331 4864 10347 4928
rect 10411 4864 10427 4928
rect 10491 4864 10507 4928
rect 10571 4864 10579 4928
rect 10259 4130 10579 4864
rect 10259 3894 10301 4130
rect 10537 3894 10579 4130
rect 10259 3840 10579 3894
rect 10259 3776 10267 3840
rect 10331 3776 10347 3840
rect 10411 3776 10427 3840
rect 10491 3776 10507 3840
rect 10571 3776 10579 3840
rect 10259 2752 10579 3776
rect 10259 2688 10267 2752
rect 10331 2688 10347 2752
rect 10411 2688 10427 2752
rect 10491 2688 10507 2752
rect 10571 2688 10579 2752
rect 10259 2128 10579 2688
rect 10919 16352 11239 16912
rect 10919 16288 10927 16352
rect 10991 16288 11007 16352
rect 11071 16288 11087 16352
rect 11151 16288 11167 16352
rect 11231 16288 11239 16352
rect 10919 15806 11239 16288
rect 10919 15570 10961 15806
rect 11197 15570 11239 15806
rect 10919 15264 11239 15570
rect 10919 15200 10927 15264
rect 10991 15200 11007 15264
rect 11071 15200 11087 15264
rect 11151 15200 11167 15264
rect 11231 15200 11239 15264
rect 10919 14176 11239 15200
rect 10919 14112 10927 14176
rect 10991 14112 11007 14176
rect 11071 14112 11087 14176
rect 11151 14112 11167 14176
rect 11231 14112 11239 14176
rect 10919 13088 11239 14112
rect 10919 13024 10927 13088
rect 10991 13024 11007 13088
rect 11071 13024 11087 13088
rect 11151 13024 11167 13088
rect 11231 13024 11239 13088
rect 10919 12134 11239 13024
rect 10919 12000 10961 12134
rect 11197 12000 11239 12134
rect 10919 11936 10927 12000
rect 11231 11936 11239 12000
rect 10919 11898 10961 11936
rect 11197 11898 11239 11936
rect 10919 10912 11239 11898
rect 10919 10848 10927 10912
rect 10991 10848 11007 10912
rect 11071 10848 11087 10912
rect 11151 10848 11167 10912
rect 11231 10848 11239 10912
rect 10919 9824 11239 10848
rect 10919 9760 10927 9824
rect 10991 9760 11007 9824
rect 11071 9760 11087 9824
rect 11151 9760 11167 9824
rect 11231 9760 11239 9824
rect 10919 8736 11239 9760
rect 10919 8672 10927 8736
rect 10991 8672 11007 8736
rect 11071 8672 11087 8736
rect 11151 8672 11167 8736
rect 11231 8672 11239 8736
rect 10919 8462 11239 8672
rect 10919 8226 10961 8462
rect 11197 8226 11239 8462
rect 10919 7648 11239 8226
rect 10919 7584 10927 7648
rect 10991 7584 11007 7648
rect 11071 7584 11087 7648
rect 11151 7584 11167 7648
rect 11231 7584 11239 7648
rect 10919 6560 11239 7584
rect 10919 6496 10927 6560
rect 10991 6496 11007 6560
rect 11071 6496 11087 6560
rect 11151 6496 11167 6560
rect 11231 6496 11239 6560
rect 10919 5472 11239 6496
rect 10919 5408 10927 5472
rect 10991 5408 11007 5472
rect 11071 5408 11087 5472
rect 11151 5408 11167 5472
rect 11231 5408 11239 5472
rect 10919 4790 11239 5408
rect 10919 4554 10961 4790
rect 11197 4554 11239 4790
rect 10919 4384 11239 4554
rect 10919 4320 10927 4384
rect 10991 4320 11007 4384
rect 11071 4320 11087 4384
rect 11151 4320 11167 4384
rect 11231 4320 11239 4384
rect 10919 3296 11239 4320
rect 10919 3232 10927 3296
rect 10991 3232 11007 3296
rect 11071 3232 11087 3296
rect 11151 3232 11167 3296
rect 11231 3232 11239 3296
rect 10919 2208 11239 3232
rect 10919 2144 10927 2208
rect 10991 2144 11007 2208
rect 11071 2144 11087 2208
rect 11151 2144 11167 2208
rect 11231 2144 11239 2208
rect 10919 2128 11239 2144
rect 13985 16896 14305 16912
rect 13985 16832 13993 16896
rect 14057 16832 14073 16896
rect 14137 16832 14153 16896
rect 14217 16832 14233 16896
rect 14297 16832 14305 16896
rect 13985 15808 14305 16832
rect 13985 15744 13993 15808
rect 14057 15744 14073 15808
rect 14137 15744 14153 15808
rect 14217 15744 14233 15808
rect 14297 15744 14305 15808
rect 13985 15146 14305 15744
rect 13985 14910 14027 15146
rect 14263 14910 14305 15146
rect 13985 14720 14305 14910
rect 13985 14656 13993 14720
rect 14057 14656 14073 14720
rect 14137 14656 14153 14720
rect 14217 14656 14233 14720
rect 14297 14656 14305 14720
rect 13985 13632 14305 14656
rect 13985 13568 13993 13632
rect 14057 13568 14073 13632
rect 14137 13568 14153 13632
rect 14217 13568 14233 13632
rect 14297 13568 14305 13632
rect 13985 12544 14305 13568
rect 13985 12480 13993 12544
rect 14057 12480 14073 12544
rect 14137 12480 14153 12544
rect 14217 12480 14233 12544
rect 14297 12480 14305 12544
rect 13985 11474 14305 12480
rect 13985 11456 14027 11474
rect 14263 11456 14305 11474
rect 13985 11392 13993 11456
rect 14297 11392 14305 11456
rect 13985 11238 14027 11392
rect 14263 11238 14305 11392
rect 13985 10368 14305 11238
rect 13985 10304 13993 10368
rect 14057 10304 14073 10368
rect 14137 10304 14153 10368
rect 14217 10304 14233 10368
rect 14297 10304 14305 10368
rect 13985 9280 14305 10304
rect 13985 9216 13993 9280
rect 14057 9216 14073 9280
rect 14137 9216 14153 9280
rect 14217 9216 14233 9280
rect 14297 9216 14305 9280
rect 13985 8192 14305 9216
rect 13985 8128 13993 8192
rect 14057 8128 14073 8192
rect 14137 8128 14153 8192
rect 14217 8128 14233 8192
rect 14297 8128 14305 8192
rect 13985 7802 14305 8128
rect 13985 7566 14027 7802
rect 14263 7566 14305 7802
rect 13985 7104 14305 7566
rect 13985 7040 13993 7104
rect 14057 7040 14073 7104
rect 14137 7040 14153 7104
rect 14217 7040 14233 7104
rect 14297 7040 14305 7104
rect 13985 6016 14305 7040
rect 13985 5952 13993 6016
rect 14057 5952 14073 6016
rect 14137 5952 14153 6016
rect 14217 5952 14233 6016
rect 14297 5952 14305 6016
rect 13985 4928 14305 5952
rect 13985 4864 13993 4928
rect 14057 4864 14073 4928
rect 14137 4864 14153 4928
rect 14217 4864 14233 4928
rect 14297 4864 14305 4928
rect 13985 4130 14305 4864
rect 13985 3894 14027 4130
rect 14263 3894 14305 4130
rect 13985 3840 14305 3894
rect 13985 3776 13993 3840
rect 14057 3776 14073 3840
rect 14137 3776 14153 3840
rect 14217 3776 14233 3840
rect 14297 3776 14305 3840
rect 13985 2752 14305 3776
rect 13985 2688 13993 2752
rect 14057 2688 14073 2752
rect 14137 2688 14153 2752
rect 14217 2688 14233 2752
rect 14297 2688 14305 2752
rect 13985 2128 14305 2688
rect 14645 16352 14965 16912
rect 14645 16288 14653 16352
rect 14717 16288 14733 16352
rect 14797 16288 14813 16352
rect 14877 16288 14893 16352
rect 14957 16288 14965 16352
rect 14645 15806 14965 16288
rect 14645 15570 14687 15806
rect 14923 15570 14965 15806
rect 14645 15264 14965 15570
rect 14645 15200 14653 15264
rect 14717 15200 14733 15264
rect 14797 15200 14813 15264
rect 14877 15200 14893 15264
rect 14957 15200 14965 15264
rect 14645 14176 14965 15200
rect 14645 14112 14653 14176
rect 14717 14112 14733 14176
rect 14797 14112 14813 14176
rect 14877 14112 14893 14176
rect 14957 14112 14965 14176
rect 14645 13088 14965 14112
rect 14645 13024 14653 13088
rect 14717 13024 14733 13088
rect 14797 13024 14813 13088
rect 14877 13024 14893 13088
rect 14957 13024 14965 13088
rect 14645 12134 14965 13024
rect 14645 12000 14687 12134
rect 14923 12000 14965 12134
rect 14645 11936 14653 12000
rect 14957 11936 14965 12000
rect 14645 11898 14687 11936
rect 14923 11898 14965 11936
rect 14645 10912 14965 11898
rect 14645 10848 14653 10912
rect 14717 10848 14733 10912
rect 14797 10848 14813 10912
rect 14877 10848 14893 10912
rect 14957 10848 14965 10912
rect 14645 9824 14965 10848
rect 14645 9760 14653 9824
rect 14717 9760 14733 9824
rect 14797 9760 14813 9824
rect 14877 9760 14893 9824
rect 14957 9760 14965 9824
rect 14645 8736 14965 9760
rect 14645 8672 14653 8736
rect 14717 8672 14733 8736
rect 14797 8672 14813 8736
rect 14877 8672 14893 8736
rect 14957 8672 14965 8736
rect 14645 8462 14965 8672
rect 14645 8226 14687 8462
rect 14923 8226 14965 8462
rect 14645 7648 14965 8226
rect 14645 7584 14653 7648
rect 14717 7584 14733 7648
rect 14797 7584 14813 7648
rect 14877 7584 14893 7648
rect 14957 7584 14965 7648
rect 14645 6560 14965 7584
rect 14645 6496 14653 6560
rect 14717 6496 14733 6560
rect 14797 6496 14813 6560
rect 14877 6496 14893 6560
rect 14957 6496 14965 6560
rect 14645 5472 14965 6496
rect 14645 5408 14653 5472
rect 14717 5408 14733 5472
rect 14797 5408 14813 5472
rect 14877 5408 14893 5472
rect 14957 5408 14965 5472
rect 14645 4790 14965 5408
rect 14645 4554 14687 4790
rect 14923 4554 14965 4790
rect 14645 4384 14965 4554
rect 14645 4320 14653 4384
rect 14717 4320 14733 4384
rect 14797 4320 14813 4384
rect 14877 4320 14893 4384
rect 14957 4320 14965 4384
rect 14645 3296 14965 4320
rect 14645 3232 14653 3296
rect 14717 3232 14733 3296
rect 14797 3232 14813 3296
rect 14877 3232 14893 3296
rect 14957 3232 14965 3296
rect 14645 2208 14965 3232
rect 14645 2144 14653 2208
rect 14717 2144 14733 2208
rect 14797 2144 14813 2208
rect 14877 2144 14893 2208
rect 14957 2144 14965 2208
rect 14645 2128 14965 2144
<< via4 >>
rect 2849 14910 3085 15146
rect 2849 11456 3085 11474
rect 2849 11392 2879 11456
rect 2879 11392 2895 11456
rect 2895 11392 2959 11456
rect 2959 11392 2975 11456
rect 2975 11392 3039 11456
rect 3039 11392 3055 11456
rect 3055 11392 3085 11456
rect 2849 11238 3085 11392
rect 2849 7566 3085 7802
rect 2849 3894 3085 4130
rect 3509 15570 3745 15806
rect 3509 12000 3745 12134
rect 3509 11936 3539 12000
rect 3539 11936 3555 12000
rect 3555 11936 3619 12000
rect 3619 11936 3635 12000
rect 3635 11936 3699 12000
rect 3699 11936 3715 12000
rect 3715 11936 3745 12000
rect 3509 11898 3745 11936
rect 3509 8226 3745 8462
rect 3509 4554 3745 4790
rect 6575 14910 6811 15146
rect 6575 11456 6811 11474
rect 6575 11392 6605 11456
rect 6605 11392 6621 11456
rect 6621 11392 6685 11456
rect 6685 11392 6701 11456
rect 6701 11392 6765 11456
rect 6765 11392 6781 11456
rect 6781 11392 6811 11456
rect 6575 11238 6811 11392
rect 6575 7566 6811 7802
rect 6575 3894 6811 4130
rect 7235 15570 7471 15806
rect 7235 12000 7471 12134
rect 7235 11936 7265 12000
rect 7265 11936 7281 12000
rect 7281 11936 7345 12000
rect 7345 11936 7361 12000
rect 7361 11936 7425 12000
rect 7425 11936 7441 12000
rect 7441 11936 7471 12000
rect 7235 11898 7471 11936
rect 7235 8226 7471 8462
rect 7235 4554 7471 4790
rect 10301 14910 10537 15146
rect 10301 11456 10537 11474
rect 10301 11392 10331 11456
rect 10331 11392 10347 11456
rect 10347 11392 10411 11456
rect 10411 11392 10427 11456
rect 10427 11392 10491 11456
rect 10491 11392 10507 11456
rect 10507 11392 10537 11456
rect 10301 11238 10537 11392
rect 10301 7566 10537 7802
rect 10301 3894 10537 4130
rect 10961 15570 11197 15806
rect 10961 12000 11197 12134
rect 10961 11936 10991 12000
rect 10991 11936 11007 12000
rect 11007 11936 11071 12000
rect 11071 11936 11087 12000
rect 11087 11936 11151 12000
rect 11151 11936 11167 12000
rect 11167 11936 11197 12000
rect 10961 11898 11197 11936
rect 10961 8226 11197 8462
rect 10961 4554 11197 4790
rect 14027 14910 14263 15146
rect 14027 11456 14263 11474
rect 14027 11392 14057 11456
rect 14057 11392 14073 11456
rect 14073 11392 14137 11456
rect 14137 11392 14153 11456
rect 14153 11392 14217 11456
rect 14217 11392 14233 11456
rect 14233 11392 14263 11456
rect 14027 11238 14263 11392
rect 14027 7566 14263 7802
rect 14027 3894 14263 4130
rect 14687 15570 14923 15806
rect 14687 12000 14923 12134
rect 14687 11936 14717 12000
rect 14717 11936 14733 12000
rect 14733 11936 14797 12000
rect 14797 11936 14813 12000
rect 14813 11936 14877 12000
rect 14877 11936 14893 12000
rect 14893 11936 14923 12000
rect 14687 11898 14923 11936
rect 14687 8226 14923 8462
rect 14687 4554 14923 4790
<< metal5 >>
rect 1056 15806 16056 15848
rect 1056 15570 3509 15806
rect 3745 15570 7235 15806
rect 7471 15570 10961 15806
rect 11197 15570 14687 15806
rect 14923 15570 16056 15806
rect 1056 15528 16056 15570
rect 1056 15146 16056 15188
rect 1056 14910 2849 15146
rect 3085 14910 6575 15146
rect 6811 14910 10301 15146
rect 10537 14910 14027 15146
rect 14263 14910 16056 15146
rect 1056 14868 16056 14910
rect 1056 12134 16056 12176
rect 1056 11898 3509 12134
rect 3745 11898 7235 12134
rect 7471 11898 10961 12134
rect 11197 11898 14687 12134
rect 14923 11898 16056 12134
rect 1056 11856 16056 11898
rect 1056 11474 16056 11516
rect 1056 11238 2849 11474
rect 3085 11238 6575 11474
rect 6811 11238 10301 11474
rect 10537 11238 14027 11474
rect 14263 11238 16056 11474
rect 1056 11196 16056 11238
rect 1056 8462 16056 8504
rect 1056 8226 3509 8462
rect 3745 8226 7235 8462
rect 7471 8226 10961 8462
rect 11197 8226 14687 8462
rect 14923 8226 16056 8462
rect 1056 8184 16056 8226
rect 1056 7802 16056 7844
rect 1056 7566 2849 7802
rect 3085 7566 6575 7802
rect 6811 7566 10301 7802
rect 10537 7566 14027 7802
rect 14263 7566 16056 7802
rect 1056 7524 16056 7566
rect 1056 4790 16056 4832
rect 1056 4554 3509 4790
rect 3745 4554 7235 4790
rect 7471 4554 10961 4790
rect 11197 4554 14687 4790
rect 14923 4554 16056 4790
rect 1056 4512 16056 4554
rect 1056 4130 16056 4172
rect 1056 3894 2849 4130
rect 3085 3894 6575 4130
rect 6811 3894 10301 4130
rect 10537 3894 14027 4130
rect 14263 3894 16056 4130
rect 1056 3852 16056 3894
use sky130_fd_sc_hd__inv_2  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1723858470
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1723858470
transform 1 0 9108 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1723858470
transform -1 0 10212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9660 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _162_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 10672 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1723858470
transform -1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 12788 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1723858470
transform -1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1723858470
transform 1 0 5152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1723858470
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3220 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1723858470
transform -1 0 4140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _171_
timestamp 1723858470
transform 1 0 3220 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1723858470
transform -1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1723858470
transform -1 0 6256 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1723858470
transform 1 0 7636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_2  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7176 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _177_
timestamp 1723858470
transform -1 0 8924 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1723858470
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1723858470
transform 1 0 13616 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _182_
timestamp 1723858470
transform 1 0 13064 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1723858470
transform 1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _185_
timestamp 1723858470
transform 1 0 14720 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _186_
timestamp 1723858470
transform -1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12328 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1723858470
transform -1 0 13984 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _189_
timestamp 1723858470
transform -1 0 12144 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _190_
timestamp 1723858470
transform -1 0 8556 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _191_
timestamp 1723858470
transform -1 0 5244 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _192_
timestamp 1723858470
transform -1 0 15180 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_2  _193_
timestamp 1723858470
transform 1 0 10764 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _194_
timestamp 1723858470
transform -1 0 6992 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _195_
timestamp 1723858470
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _196_
timestamp 1723858470
transform -1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _197_
timestamp 1723858470
transform -1 0 13984 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _198_
timestamp 1723858470
transform -1 0 11408 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6716 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _200_
timestamp 1723858470
transform 1 0 4048 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _201_
timestamp 1723858470
transform -1 0 4416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp 1723858470
transform -1 0 13616 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _203_
timestamp 1723858470
transform -1 0 12236 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _204_
timestamp 1723858470
transform -1 0 8464 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _205_
timestamp 1723858470
transform 1 0 5060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _206_
timestamp 1723858470
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _207_
timestamp 1723858470
transform -1 0 4876 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _208_
timestamp 1723858470
transform -1 0 13340 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _210_
timestamp 1723858470
transform -1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7636 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _214_
timestamp 1723858470
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _215_
timestamp 1723858470
transform -1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _216_
timestamp 1723858470
transform -1 0 5520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _217_
timestamp 1723858470
transform -1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _218_
timestamp 1723858470
transform -1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _219_
timestamp 1723858470
transform -1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _220_
timestamp 1723858470
transform -1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5244 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _223_
timestamp 1723858470
transform 1 0 7084 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _224_
timestamp 1723858470
transform 1 0 5060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6256 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _227_
timestamp 1723858470
transform -1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _228_
timestamp 1723858470
transform 1 0 4600 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _229_
timestamp 1723858470
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4048 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _231_
timestamp 1723858470
transform -1 0 3128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _232_
timestamp 1723858470
transform -1 0 5520 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _233_
timestamp 1723858470
transform -1 0 5152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _235_
timestamp 1723858470
transform -1 0 4784 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _236_
timestamp 1723858470
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4968 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _238_
timestamp 1723858470
transform 1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _239_
timestamp 1723858470
transform -1 0 3496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _240_
timestamp 1723858470
transform -1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _241_
timestamp 1723858470
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp 1723858470
transform -1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _243_
timestamp 1723858470
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8096 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _245_
timestamp 1723858470
transform -1 0 8740 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _246_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 11316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _247_
timestamp 1723858470
transform 1 0 9108 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6716 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _249_
timestamp 1723858470
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _250_
timestamp 1723858470
transform 1 0 2392 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _251_
timestamp 1723858470
transform 1 0 7544 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8740 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _253_
timestamp 1723858470
transform -1 0 9568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _254_
timestamp 1723858470
transform 1 0 9660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _255_
timestamp 1723858470
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _256_
timestamp 1723858470
transform 1 0 7820 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _257_
timestamp 1723858470
transform -1 0 6164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _258_
timestamp 1723858470
transform 1 0 7728 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _260_
timestamp 1723858470
transform -1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _261_
timestamp 1723858470
transform 1 0 7728 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _262_
timestamp 1723858470
transform 1 0 5612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp 1723858470
transform 1 0 4784 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _264_
timestamp 1723858470
transform 1 0 8188 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _265_
timestamp 1723858470
transform 1 0 7820 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _266_
timestamp 1723858470
transform 1 0 5060 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _267_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6532 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7176 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _269_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 12328 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _271_
timestamp 1723858470
transform -1 0 12788 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _272_
timestamp 1723858470
transform 1 0 12328 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _273_
timestamp 1723858470
transform -1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _274_
timestamp 1723858470
transform -1 0 13708 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _275_
timestamp 1723858470
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _276_
timestamp 1723858470
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1723858470
transform 1 0 10120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _278_
timestamp 1723858470
transform 1 0 3864 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 12604 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _280_
timestamp 1723858470
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _281_
timestamp 1723858470
transform 1 0 12604 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1723858470
transform -1 0 12512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _283_
timestamp 1723858470
transform -1 0 12880 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _284_
timestamp 1723858470
transform 1 0 11592 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _285_
timestamp 1723858470
transform 1 0 10212 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _286_
timestamp 1723858470
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _287_
timestamp 1723858470
transform -1 0 13984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _288_
timestamp 1723858470
transform -1 0 11224 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _289_
timestamp 1723858470
transform 1 0 10672 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _290_
timestamp 1723858470
transform 1 0 10764 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _291_
timestamp 1723858470
transform -1 0 10856 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _292_
timestamp 1723858470
transform 1 0 10856 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _293_
timestamp 1723858470
transform 1 0 10948 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _294_
timestamp 1723858470
transform 1 0 9660 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _295_
timestamp 1723858470
transform 1 0 11592 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _296_
timestamp 1723858470
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _297_
timestamp 1723858470
transform 1 0 9200 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 14628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _299_
timestamp 1723858470
transform 1 0 14812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _300_
timestamp 1723858470
transform -1 0 14720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _301_
timestamp 1723858470
transform -1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _302_
timestamp 1723858470
transform -1 0 8832 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _303_
timestamp 1723858470
transform 1 0 8280 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _304_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 14076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _305_
timestamp 1723858470
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _306_
timestamp 1723858470
transform 1 0 14812 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _307_
timestamp 1723858470
transform 1 0 14904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _308_
timestamp 1723858470
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _309_
timestamp 1723858470
transform -1 0 13616 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _310_
timestamp 1723858470
transform 1 0 14076 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _311_
timestamp 1723858470
transform 1 0 13156 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _312_
timestamp 1723858470
transform -1 0 15088 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _313_
timestamp 1723858470
transform 1 0 14812 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _314_
timestamp 1723858470
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _315_
timestamp 1723858470
transform 1 0 13156 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _316_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 11960 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _317_
timestamp 1723858470
transform 1 0 1840 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _318_
timestamp 1723858470
transform 1 0 4232 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _319_
timestamp 1723858470
transform 1 0 1840 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 1723858470
transform 1 0 1840 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 1723858470
transform 1 0 6348 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1723858470
transform 1 0 2760 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _323_
timestamp 1723858470
transform 1 0 1840 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _324_
timestamp 1723858470
transform 1 0 1840 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _325_
timestamp 1723858470
transform 1 0 4416 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1723858470
transform 1 0 1840 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _327_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2116 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _328_
timestamp 1723858470
transform 1 0 1748 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _329_
timestamp 1723858470
transform 1 0 1840 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _330_
timestamp 1723858470
transform 1 0 1932 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _331_
timestamp 1723858470
transform 1 0 6164 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _332_
timestamp 1723858470
transform 1 0 8924 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _333_
timestamp 1723858470
transform 1 0 6532 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _334_
timestamp 1723858470
transform 1 0 1840 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _335_
timestamp 1723858470
transform 1 0 6440 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _336_
timestamp 1723858470
transform 1 0 8924 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _337_
timestamp 1723858470
transform 1 0 6900 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _338_
timestamp 1723858470
transform 1 0 6348 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _339_
timestamp 1723858470
transform 1 0 6440 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _340_
timestamp 1723858470
transform 1 0 6992 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _341_
timestamp 1723858470
transform 1 0 4416 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _342_
timestamp 1723858470
transform 1 0 6256 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _343_
timestamp 1723858470
transform 1 0 4600 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _344_
timestamp 1723858470
transform -1 0 8280 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _345_
timestamp 1723858470
transform 1 0 5152 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _346_
timestamp 1723858470
transform 1 0 9936 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _347_
timestamp 1723858470
transform 1 0 12972 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _348_
timestamp 1723858470
transform 1 0 9568 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _349_
timestamp 1723858470
transform 1 0 3220 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _350_
timestamp 1723858470
transform 1 0 10212 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _351_
timestamp 1723858470
transform 1 0 12696 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _352_
timestamp 1723858470
transform 1 0 9752 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _353_
timestamp 1723858470
transform 1 0 9476 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _354_
timestamp 1723858470
transform 1 0 9660 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _355_
timestamp 1723858470
transform 1 0 11316 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _356_
timestamp 1723858470
transform 1 0 9108 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _357_
timestamp 1723858470
transform 1 0 9568 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _358_
timestamp 1723858470
transform 1 0 9384 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _359_
timestamp 1723858470
transform 1 0 11500 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _360_
timestamp 1723858470
transform 1 0 8832 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _361_
timestamp 1723858470
transform 1 0 13064 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _362_
timestamp 1723858470
transform 1 0 13524 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _363_
timestamp 1723858470
transform 1 0 7912 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _364_
timestamp 1723858470
transform 1 0 12144 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _365_
timestamp 1723858470
transform 1 0 13340 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _366_
timestamp 1723858470
transform 1 0 12144 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _367_
timestamp 1723858470
transform -1 0 14996 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _368_
timestamp 1723858470
transform 1 0 13708 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _369_
timestamp 1723858470
transform -1 0 14812 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _370_
timestamp 1723858470
transform -1 0 15640 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _371_
timestamp 1723858470
transform 1 0 12788 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8740 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1723858470
transform -1 0 6256 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1723858470
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1723858470
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1723858470
transform 1 0 9568 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  fanout6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9200 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 9292 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout8
timestamp 1723858470
transform -1 0 15548 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout9
timestamp 1723858470
transform -1 0 15364 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1723858470
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1723858470
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1723858470
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1723858470
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1723858470
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1723858470
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1723858470
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_100
timestamp 1723858470
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1723858470
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_125 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 1723858470
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1723858470
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_141 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_153
timestamp 1723858470
transform 1 0 15180 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1723858470
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_15
timestamp 1723858470
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1723858470
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1723858470
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1723858470
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1723858470
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1723858470
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_76
timestamp 1723858470
transform 1 0 8096 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_88
timestamp 1723858470
transform 1 0 9200 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_96
timestamp 1723858470
transform 1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 1723858470
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_113
timestamp 1723858470
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_121
timestamp 1723858470
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_156
timestamp 1723858470
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3
timestamp 1723858470
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_7
timestamp 1723858470
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_37
timestamp 1723858470
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_76
timestamp 1723858470
transform 1 0 8096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1723858470
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_85
timestamp 1723858470
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_91
timestamp 1723858470
transform 1 0 9476 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_95
timestamp 1723858470
transform 1 0 9844 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_119
timestamp 1723858470
transform 1 0 12052 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_157
timestamp 1723858470
transform 1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_3
timestamp 1723858470
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_7
timestamp 1723858470
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1723858470
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_78
timestamp 1723858470
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_88
timestamp 1723858470
transform 1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1723858470
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_158
timestamp 1723858470
transform 1 0 15640 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_3
timestamp 1723858470
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_7
timestamp 1723858470
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_56
timestamp 1723858470
transform 1 0 6256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1723858470
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1723858470
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_15
timestamp 1723858470
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_40
timestamp 1723858470
transform 1 0 4784 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_52
timestamp 1723858470
transform 1 0 5888 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_64
timestamp 1723858470
transform 1 0 6992 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_75
timestamp 1723858470
transform 1 0 8004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_87
timestamp 1723858470
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_96
timestamp 1723858470
transform 1 0 9936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1723858470
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_131
timestamp 1723858470
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_155
timestamp 1723858470
transform 1 0 15364 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1723858470
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_15
timestamp 1723858470
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1723858470
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_33
timestamp 1723858470
transform 1 0 4140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_45
timestamp 1723858470
transform 1 0 5244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_57
timestamp 1723858470
transform 1 0 6348 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_66
timestamp 1723858470
transform 1 0 7176 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_78
timestamp 1723858470
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1723858470
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_97
timestamp 1723858470
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_125
timestamp 1723858470
transform 1 0 12604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_137
timestamp 1723858470
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_148
timestamp 1723858470
transform 1 0 14720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_157
timestamp 1723858470
transform 1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1723858470
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_15
timestamp 1723858470
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_45
timestamp 1723858470
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_53
timestamp 1723858470
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1723858470
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_65
timestamp 1723858470
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1723858470
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_81
timestamp 1723858470
transform 1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_89
timestamp 1723858470
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_121
timestamp 1723858470
transform 1 0 12236 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_133
timestamp 1723858470
transform 1 0 13340 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_145
timestamp 1723858470
transform 1 0 14444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_157
timestamp 1723858470
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1723858470
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_7
timestamp 1723858470
transform 1 0 1748 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 1723858470
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_56
timestamp 1723858470
transform 1 0 6256 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_60
timestamp 1723858470
transform 1 0 6624 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1723858470
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1723858470
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1723858470
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_97
timestamp 1723858470
transform 1 0 10028 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_128
timestamp 1723858470
transform 1 0 12880 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_147
timestamp 1723858470
transform 1 0 14628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_152
timestamp 1723858470
transform 1 0 15088 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_158
timestamp 1723858470
transform 1 0 15640 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1723858470
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_41
timestamp 1723858470
transform 1 0 4876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 1723858470
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_96
timestamp 1723858470
transform 1 0 9936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_108
timestamp 1723858470
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_116
timestamp 1723858470
transform 1 0 11776 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1723858470
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_15
timestamp 1723858470
transform 1 0 2484 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_23
timestamp 1723858470
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_29
timestamp 1723858470
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_112
timestamp 1723858470
transform 1 0 11408 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_157
timestamp 1723858470
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1723858470
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_15
timestamp 1723858470
transform 1 0 2484 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_44
timestamp 1723858470
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_88
timestamp 1723858470
transform 1 0 9200 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_124
timestamp 1723858470
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_157
timestamp 1723858470
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 1723858470
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_7
timestamp 1723858470
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1723858470
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_39
timestamp 1723858470
transform 1 0 4692 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_49
timestamp 1723858470
transform 1 0 5612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_61
timestamp 1723858470
transform 1 0 6716 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1723858470
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_115
timestamp 1723858470
transform 1 0 11684 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_152
timestamp 1723858470
transform 1 0 15088 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1723858470
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_15
timestamp 1723858470
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 1723858470
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1723858470
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1723858470
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_81
timestamp 1723858470
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_103
timestamp 1723858470
transform 1 0 10580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1723858470
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1723858470
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_120
timestamp 1723858470
transform 1 0 12144 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_132
timestamp 1723858470
transform 1 0 13248 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_153
timestamp 1723858470
transform 1 0 15180 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1723858470
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_15
timestamp 1723858470
transform 1 0 2484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1723858470
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1723858470
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_41
timestamp 1723858470
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1723858470
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1723858470
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_93
timestamp 1723858470
transform 1 0 9660 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_114
timestamp 1723858470
transform 1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_125
timestamp 1723858470
transform 1 0 12604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1723858470
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_156
timestamp 1723858470
transform 1 0 15456 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_6
timestamp 1723858470
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_37
timestamp 1723858470
transform 1 0 4508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_45
timestamp 1723858470
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1723858470
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_57
timestamp 1723858470
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_89
timestamp 1723858470
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_124
timestamp 1723858470
transform 1 0 12512 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_130
timestamp 1723858470
transform 1 0 13064 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1723858470
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_15
timestamp 1723858470
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_65
timestamp 1723858470
transform 1 0 7084 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_71
timestamp 1723858470
transform 1 0 7636 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 1723858470
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_113
timestamp 1723858470
transform 1 0 11500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_128
timestamp 1723858470
transform 1 0 12880 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_155
timestamp 1723858470
transform 1 0 15364 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1723858470
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_11
timestamp 1723858470
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_20
timestamp 1723858470
transform 1 0 2944 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1723858470
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_85
timestamp 1723858470
transform 1 0 8924 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_93
timestamp 1723858470
transform 1 0 9660 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_99
timestamp 1723858470
transform 1 0 10212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1723858470
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_120
timestamp 1723858470
transform 1 0 12144 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_126
timestamp 1723858470
transform 1 0 12696 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_148
timestamp 1723858470
transform 1 0 14720 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_156
timestamp 1723858470
transform 1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_3
timestamp 1723858470
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_7
timestamp 1723858470
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_29
timestamp 1723858470
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_47
timestamp 1723858470
transform 1 0 5428 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_56
timestamp 1723858470
transform 1 0 6256 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 1723858470
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1723858470
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_104
timestamp 1723858470
transform 1 0 10672 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1723858470
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1723858470
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_150
timestamp 1723858470
transform 1 0 14904 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_158
timestamp 1723858470
transform 1 0 15640 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1723858470
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_7
timestamp 1723858470
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_29
timestamp 1723858470
transform 1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_42
timestamp 1723858470
transform 1 0 4968 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1723858470
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_69
timestamp 1723858470
transform 1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_82
timestamp 1723858470
transform 1 0 8648 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1723858470
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp 1723858470
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_119
timestamp 1723858470
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_128
timestamp 1723858470
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_140
timestamp 1723858470
transform 1 0 13984 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_152
timestamp 1723858470
transform 1 0 15088 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_158
timestamp 1723858470
transform 1 0 15640 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_3
timestamp 1723858470
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_37
timestamp 1723858470
transform 1 0 4508 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_49
timestamp 1723858470
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_61
timestamp 1723858470
transform 1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_85
timestamp 1723858470
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_96
timestamp 1723858470
transform 1 0 9936 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_112
timestamp 1723858470
transform 1 0 11408 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_124
timestamp 1723858470
transform 1 0 12512 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_130
timestamp 1723858470
transform 1 0 13064 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1723858470
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_148
timestamp 1723858470
transform 1 0 14720 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_156
timestamp 1723858470
transform 1 0 15456 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1723858470
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_21
timestamp 1723858470
transform 1 0 3036 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_32
timestamp 1723858470
transform 1 0 4048 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_40
timestamp 1723858470
transform 1 0 4784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_49
timestamp 1723858470
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1723858470
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1723858470
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1723858470
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_81
timestamp 1723858470
transform 1 0 8556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_85
timestamp 1723858470
transform 1 0 8924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_101
timestamp 1723858470
transform 1 0 10396 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1723858470
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1723858470
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_125
timestamp 1723858470
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_157
timestamp 1723858470
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1723858470
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1723858470
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1723858470
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_29
timestamp 1723858470
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_37
timestamp 1723858470
transform 1 0 4508 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_80
timestamp 1723858470
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1723858470
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_110
timestamp 1723858470
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_129
timestamp 1723858470
transform 1 0 12972 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1723858470
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_157
timestamp 1723858470
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1723858470
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_15
timestamp 1723858470
transform 1 0 2484 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_21
timestamp 1723858470
transform 1 0 3036 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_26
timestamp 1723858470
transform 1 0 3496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1723858470
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_84
timestamp 1723858470
transform 1 0 8832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1723858470
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1723858470
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_117
timestamp 1723858470
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_158
timestamp 1723858470
transform 1 0 15640 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 1723858470
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_7
timestamp 1723858470
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_37
timestamp 1723858470
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1723858470
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_85
timestamp 1723858470
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_100
timestamp 1723858470
transform 1 0 10304 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_112
timestamp 1723858470
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 1723858470
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1723858470
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_153
timestamp 1723858470
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1723858470
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_15
timestamp 1723858470
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1723858470
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1723858470
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_57
timestamp 1723858470
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_63
timestamp 1723858470
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_72
timestamp 1723858470
transform 1 0 7728 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_95
timestamp 1723858470
transform 1 0 9844 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_103
timestamp 1723858470
transform 1 0 10580 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_121
timestamp 1723858470
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_130
timestamp 1723858470
transform 1 0 13064 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_142
timestamp 1723858470
transform 1 0 14168 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_154
timestamp 1723858470
transform 1 0 15272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_158
timestamp 1723858470
transform 1 0 15640 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1723858470
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1723858470
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1723858470
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_29
timestamp 1723858470
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_37
timestamp 1723858470
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_48
timestamp 1723858470
transform 1 0 5520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_57
timestamp 1723858470
transform 1 0 6348 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_65
timestamp 1723858470
transform 1 0 7084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 1723858470
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1723858470
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1723858470
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_109
timestamp 1723858470
transform 1 0 11132 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_113
timestamp 1723858470
transform 1 0 11500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1723858470
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1723858470
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1723858470
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1723858470
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_153
timestamp 1723858470
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 15548 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1723858470
transform 1 0 12972 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1723858470
transform -1 0 12880 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1723858470
transform -1 0 6256 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1723858470
transform -1 0 13064 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1723858470
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1723858470
transform -1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1723858470
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1723858470
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1723858470
transform -1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8464 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1723858470
transform 1 0 3956 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1723858470
transform 1 0 3772 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1723858470
transform -1 0 6256 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1723858470
transform -1 0 5428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1723858470
transform -1 0 10764 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1723858470
transform -1 0 9936 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1723858470
transform -1 0 8004 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1723858470
transform -1 0 5796 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1723858470
transform -1 0 7176 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1723858470
transform -1 0 4048 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1723858470
transform 1 0 14996 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1723858470
transform -1 0 14812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1723858470
transform -1 0 12880 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1723858470
transform -1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1723858470
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1723858470
transform -1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1723858470
transform -1 0 5520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1723858470
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1723858470
transform -1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1723858470
transform -1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1723858470
transform -1 0 10672 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1723858470
transform -1 0 9936 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1723858470
transform 1 0 11868 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1723858470
transform -1 0 9660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1723858470
transform -1 0 7636 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1723858470
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1723858470
transform -1 0 10948 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1723858470
transform -1 0 14904 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1723858470
transform -1 0 11408 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1723858470
transform -1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1723858470
transform -1 0 9108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1723858470
transform -1 0 12328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1723858470
transform -1 0 3772 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1723858470
transform 1 0 12328 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1723858470
transform 1 0 3956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1723858470
transform -1 0 8556 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1723858470
transform 1 0 6992 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1723858470
transform 1 0 11776 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1723858470
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1723858470
transform 1 0 3864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1723858470
transform 1 0 14812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1723858470
transform -1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1723858470
transform -1 0 4508 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1723858470
transform 1 0 4140 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1723858470
transform -1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1723858470
transform -1 0 7176 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1723858470
transform -1 0 15732 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1723858470
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1723858470
transform 1 0 9752 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1723858470
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1723858470
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1723858470
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1723858470
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1723858470
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1723858470
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1723858470
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1723858470
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1723858470
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1723858470
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1723858470
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1723858470
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1723858470
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1723858470
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1723858470
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1723858470
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1723858470
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1723858470
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1723858470
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1723858470
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1723858470
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1723858470
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1723858470
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1723858470
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1723858470
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1723858470
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1723858470
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1723858470
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1723858470
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1723858470
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1723858470
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1723858470
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1723858470
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1723858470
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1723858470
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1723858470
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1723858470
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1723858470
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1723858470
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1723858470
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1723858470
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1723858470
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1723858470
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1723858470
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1723858470
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1723858470
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1723858470
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1723858470
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1723858470
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1723858470
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1723858470
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1723858470
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1723858470
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1723858470
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1723858470
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1723858470
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1723858470
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1723858470
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1723858470
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1723858470
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1723858470
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1723858470
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1723858470
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1723858470
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1723858470
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1723858470
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1723858470
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1723858470
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1723858470
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1723858470
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1723858470
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1723858470
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1723858470
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1723858470
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1723858470
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1723858470
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1723858470
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1723858470
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1723858470
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1723858470
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1723858470
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1723858470
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1723858470
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1723858470
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1723858470
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1723858470
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1723858470
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1723858470
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1723858470
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1723858470
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1723858470
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1723858470
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1723858470
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1723858470
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1723858470
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1723858470
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1723858470
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1723858470
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1723858470
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1723858470
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1723858470
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1723858470
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1723858470
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1723858470
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1723858470
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1723858470
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1723858470
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1723858470
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1723858470
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1723858470
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1723858470
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1723858470
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1723858470
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1723858470
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1723858470
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1723858470
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1723858470
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1723858470
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1723858470
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1723858470
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1723858470
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1723858470
transform 1 0 6256 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1723858470
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1723858470
transform 1 0 11408 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1723858470
transform 1 0 13984 0 1 16320
box -38 -48 130 592
<< labels >>
flabel metal4 s 3467 2128 3787 16912 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7193 2128 7513 16912 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10919 2128 11239 16912 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14645 2128 14965 16912 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4512 16056 4832 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8184 16056 8504 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 11856 16056 12176 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 15528 16056 15848 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2807 2128 3127 16912 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6533 2128 6853 16912 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 10259 2128 10579 16912 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13985 2128 14305 16912 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3852 16056 4172 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7524 16056 7844 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 11196 16056 11516 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 14868 16056 15188 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 13542 18546 13598 19346 0 FreeSans 224 90 0 0 a_in[0]
port 2 nsew signal input
flabel metal2 s 7102 18546 7158 19346 0 FreeSans 224 90 0 0 a_in[1]
port 3 nsew signal input
flabel metal3 s 16402 15648 17202 15768 0 FreeSans 480 0 0 0 a_in[2]
port 4 nsew signal input
flabel metal3 s 16402 5448 17202 5568 0 FreeSans 480 0 0 0 a_in[3]
port 5 nsew signal input
flabel metal2 s 3882 18546 3938 19346 0 FreeSans 224 90 0 0 a_in[4]
port 6 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 a_in[5]
port 7 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 a_in[6]
port 8 nsew signal input
flabel metal3 s 16402 2048 17202 2168 0 FreeSans 480 0 0 0 a_in[7]
port 9 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 a_in_ready
port 10 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 a_in_valid
port 11 nsew signal input
flabel metal2 s 16762 18546 16818 19346 0 FreeSans 224 90 0 0 b_in[0]
port 12 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 b_in[1]
port 13 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 b_in[2]
port 14 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 b_in[3]
port 15 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 b_in[4]
port 16 nsew signal input
flabel metal3 s 16402 12248 17202 12368 0 FreeSans 480 0 0 0 b_in[5]
port 17 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 b_in[6]
port 18 nsew signal input
flabel metal2 s 10322 18546 10378 19346 0 FreeSans 224 90 0 0 b_in[7]
port 19 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 b_in_ready
port 20 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 b_in_valid
port 21 nsew signal input
flabel metal2 s 662 18546 718 19346 0 FreeSans 224 90 0 0 clk
port 22 nsew signal input
flabel metal3 s 16402 8848 17202 8968 0 FreeSans 480 0 0 0 rst_n
port 23 nsew signal input
rlabel metal1 8556 16320 8556 16320 0 VGND
rlabel metal1 8556 16864 8556 16864 0 VPWR
rlabel metal2 12282 14756 12282 14756 0 _000_
rlabel metal2 2162 3298 2162 3298 0 _001_
rlabel metal1 4738 3706 4738 3706 0 _002_
rlabel metal1 2346 4658 2346 4658 0 _003_
rlabel metal1 4692 6426 4692 6426 0 _004_
rlabel metal1 6164 6630 6164 6630 0 _005_
rlabel metal1 3864 8398 3864 8398 0 _006_
rlabel metal2 3174 4794 3174 4794 0 _007_
rlabel metal1 4094 9078 4094 9078 0 _008_
rlabel metal1 5106 11322 5106 11322 0 _009_
rlabel metal1 2162 12104 2162 12104 0 _010_
rlabel metal2 4922 7106 4922 7106 0 _011_
rlabel metal1 2300 13362 2300 13362 0 _012_
rlabel metal1 2162 15368 2162 15368 0 _013_
rlabel metal2 2254 10404 2254 10404 0 _014_
rlabel metal1 7590 3570 7590 3570 0 _015_
rlabel metal1 9614 3706 9614 3706 0 _016_
rlabel metal1 7636 4658 7636 4658 0 _017_
rlabel metal1 2300 11866 2300 11866 0 _018_
rlabel metal1 7406 6970 7406 6970 0 _019_
rlabel metal1 9476 7922 9476 7922 0 _020_
rlabel metal1 7544 10234 7544 10234 0 _021_
rlabel metal2 6118 3808 6118 3808 0 _022_
rlabel metal1 7682 11322 7682 11322 0 _023_
rlabel metal1 7682 12954 7682 12954 0 _024_
rlabel metal1 4784 14586 4784 14586 0 _025_
rlabel metal1 8142 8058 8142 8058 0 _026_
rlabel metal1 5336 14518 5336 14518 0 _027_
rlabel metal1 7130 16150 7130 16150 0 _028_
rlabel metal1 5513 11322 5513 11322 0 _029_
rlabel metal1 10987 3706 10987 3706 0 _030_
rlabel metal1 13524 4046 13524 4046 0 _031_
rlabel metal1 10028 5882 10028 5882 0 _032_
rlabel metal2 3910 15572 3910 15572 0 _033_
rlabel metal2 11546 6698 11546 6698 0 _034_
rlabel metal1 12742 8534 12742 8534 0 _035_
rlabel metal1 11500 9622 11500 9622 0 _036_
rlabel metal1 10028 3162 10028 3162 0 _037_
rlabel metal1 11454 10778 11454 10778 0 _038_
rlabel metal1 11638 12104 11638 12104 0 _039_
rlabel metal2 11086 13668 11086 13668 0 _040_
rlabel metal1 10948 9010 10948 9010 0 _041_
rlabel metal2 9706 15198 9706 15198 0 _042_
rlabel metal1 11316 16014 11316 16014 0 _043_
rlabel metal1 9522 12342 9522 12342 0 _044_
rlabel metal1 13386 3128 13386 3128 0 _045_
rlabel metal1 13984 5270 13984 5270 0 _046_
rlabel metal1 8280 15674 8280 15674 0 _047_
rlabel metal1 13984 6970 13984 6970 0 _048_
rlabel metal1 13800 9622 13800 9622 0 _049_
rlabel metal1 14996 3094 14996 3094 0 _050_
rlabel metal1 14628 10710 14628 10710 0 _051_
rlabel metal1 13248 13498 13248 13498 0 _052_
rlabel metal1 15042 7446 15042 7446 0 _053_
rlabel metal1 15042 14586 15042 14586 0 _054_
rlabel metal1 13156 11798 13156 11798 0 _055_
rlabel metal2 11546 4896 11546 4896 0 _056_
rlabel metal1 11408 9486 11408 9486 0 _057_
rlabel metal1 9430 13940 9430 13940 0 _058_
rlabel metal1 8602 12852 8602 12852 0 _059_
rlabel metal1 9262 12206 9262 12206 0 _060_
rlabel metal1 11960 8942 11960 8942 0 _061_
rlabel metal2 12834 4998 12834 4998 0 _062_
rlabel metal2 12558 4573 12558 4573 0 _063_
rlabel metal1 4370 4556 4370 4556 0 _064_
rlabel metal1 3910 9588 3910 9588 0 _065_
rlabel metal1 3818 9520 3818 9520 0 _066_
rlabel metal1 3312 9554 3312 9554 0 _067_
rlabel metal1 3450 6222 3450 6222 0 _068_
rlabel metal1 4048 6902 4048 6902 0 _069_
rlabel metal1 3910 4046 3910 4046 0 _070_
rlabel metal1 4738 4794 4738 4794 0 _071_
rlabel metal1 11592 4114 11592 4114 0 _072_
rlabel metal1 6394 5236 6394 5236 0 _073_
rlabel metal1 7314 12138 7314 12138 0 _074_
rlabel metal1 7176 14246 7176 14246 0 _075_
rlabel metal1 8648 9078 8648 9078 0 _076_
rlabel metal1 7774 5236 7774 5236 0 _077_
rlabel metal1 11500 4182 11500 4182 0 _078_
rlabel metal2 15502 4386 15502 4386 0 _079_
rlabel metal1 13064 14382 13064 14382 0 _080_
rlabel metal1 13478 12614 13478 12614 0 _081_
rlabel metal1 14858 8908 14858 8908 0 _082_
rlabel metal1 14214 6630 14214 6630 0 _083_
rlabel metal1 14306 6800 14306 6800 0 _084_
rlabel metal1 12466 4182 12466 4182 0 _085_
rlabel metal1 13616 12818 13616 12818 0 _086_
rlabel metal2 8556 12580 8556 12580 0 _087_
rlabel metal2 5244 12716 5244 12716 0 _088_
rlabel metal1 4232 9690 4232 9690 0 _089_
rlabel metal2 13202 3536 13202 3536 0 _090_
rlabel metal2 10994 4828 10994 4828 0 _091_
rlabel metal1 5428 3502 5428 3502 0 _092_
rlabel metal1 4232 4794 4232 4794 0 _093_
rlabel metal1 11822 7922 11822 7922 0 _094_
rlabel metal1 12374 9010 12374 9010 0 _095_
rlabel metal1 7268 8942 7268 8942 0 _096_
rlabel metal1 5612 7514 5612 7514 0 _097_
rlabel metal1 4416 7514 4416 7514 0 _098_
rlabel metal2 4278 11492 4278 11492 0 _099_
rlabel metal2 13386 14501 13386 14501 0 _100_
rlabel metal2 9890 15028 9890 15028 0 _101_
rlabel metal1 6486 14926 6486 14926 0 _102_
rlabel metal1 4784 14042 4784 14042 0 _103_
rlabel metal1 4554 7412 4554 7412 0 _104_
rlabel metal1 13018 14246 13018 14246 0 _105_
rlabel metal2 2714 4896 2714 4896 0 _106_
rlabel metal1 6624 4998 6624 4998 0 _107_
rlabel metal2 2714 10387 2714 10387 0 _108_
rlabel metal2 3910 6171 3910 6171 0 _109_
rlabel metal1 4968 4658 4968 4658 0 _110_
rlabel metal1 5244 4794 5244 4794 0 _111_
rlabel metal1 5060 3570 5060 3570 0 _112_
rlabel metal1 3588 4046 3588 4046 0 _113_
rlabel metal1 5382 6970 5382 6970 0 _114_
rlabel metal1 7866 6800 7866 6800 0 _115_
rlabel metal1 5060 7242 5060 7242 0 _116_
rlabel metal1 6118 6766 6118 6766 0 _117_
rlabel metal1 4876 8466 4876 8466 0 _118_
rlabel metal1 4646 11084 4646 11084 0 _119_
rlabel metal1 5106 12954 5106 12954 0 _120_
rlabel metal1 4416 11186 4416 11186 0 _121_
rlabel metal1 2668 11730 2668 11730 0 _122_
rlabel metal1 3036 14926 3036 14926 0 _123_
rlabel metal2 8418 7684 8418 7684 0 _124_
rlabel metal1 6946 5712 6946 5712 0 _125_
rlabel metal1 7314 3060 7314 3060 0 _126_
rlabel metal1 9430 3604 9430 3604 0 _127_
rlabel metal1 8372 4590 8372 4590 0 _128_
rlabel metal1 9108 9146 9108 9146 0 _129_
rlabel metal1 9522 8602 9522 8602 0 _130_
rlabel metal1 8050 10064 8050 10064 0 _131_
rlabel metal1 5750 12784 5750 12784 0 _132_
rlabel metal1 7958 12852 7958 12852 0 _133_
rlabel metal1 5014 14416 5014 14416 0 _134_
rlabel metal1 5290 14314 5290 14314 0 _135_
rlabel metal1 7452 15130 7452 15130 0 _136_
rlabel metal1 12558 4080 12558 4080 0 _137_
rlabel metal2 12650 3638 12650 3638 0 _138_
rlabel metal1 12650 5270 12650 5270 0 _139_
rlabel metal1 13800 4590 13800 4590 0 _140_
rlabel metal2 11546 5474 11546 5474 0 _141_
rlabel metal1 12006 8874 12006 8874 0 _142_
rlabel metal2 12650 8636 12650 8636 0 _143_
rlabel metal2 12558 10234 12558 10234 0 _144_
rlabel metal1 13110 12104 13110 12104 0 _145_
rlabel metal1 11362 13362 11362 13362 0 _146_
rlabel metal2 10718 12517 10718 12517 0 _147_
rlabel metal1 10856 13362 10856 13362 0 _148_
rlabel metal1 10902 16116 10902 16116 0 _149_
rlabel metal1 14030 4794 14030 4794 0 _150_
rlabel metal1 14352 5746 14352 5746 0 _151_
rlabel metal1 8648 15130 8648 15130 0 _152_
rlabel metal1 14904 9146 14904 9146 0 _153_
rlabel metal1 13800 14314 13800 14314 0 _154_
rlabel metal1 13662 13362 13662 13362 0 _155_
rlabel metal2 15042 8092 15042 8092 0 _156_
rlabel metal2 12926 1520 12926 1520 0 a_in_ready
rlabel metal2 46 1554 46 1554 0 a_in_valid
rlabel metal2 9706 1520 9706 1520 0 b_in_ready
rlabel metal3 820 10268 820 10268 0 b_in_valid
rlabel metal2 690 14069 690 14069 0 clk
rlabel metal1 10442 9350 10442 9350 0 clknet_0_clk
rlabel metal2 1886 5746 1886 5746 0 clknet_2_0__leaf_clk
rlabel metal2 1978 11084 1978 11084 0 clknet_2_1__leaf_clk
rlabel via1 13018 3570 13018 3570 0 clknet_2_2__leaf_clk
rlabel metal1 13754 13974 13754 13974 0 clknet_2_3__leaf_clk
rlabel metal1 13570 3910 13570 3910 0 net1
rlabel metal1 14398 14246 14398 14246 0 net10
rlabel metal1 13846 13838 13846 13838 0 net11
rlabel metal2 12190 12512 12190 12512 0 net12
rlabel metal1 5658 3706 5658 3706 0 net13
rlabel metal1 11822 16150 11822 16150 0 net14
rlabel metal1 12006 15538 12006 15538 0 net15
rlabel metal2 14490 6222 14490 6222 0 net16
rlabel metal2 4278 15164 4278 15164 0 net17
rlabel metal1 11316 14042 11316 14042 0 net18
rlabel metal1 9568 14042 9568 14042 0 net19
rlabel metal1 3634 10030 3634 10030 0 net2
rlabel metal2 8602 4250 8602 4250 0 net20
rlabel metal1 3772 13906 3772 13906 0 net21
rlabel metal1 4554 5338 4554 5338 0 net22
rlabel metal1 5198 12886 5198 12886 0 net23
rlabel metal2 4738 11866 4738 11866 0 net24
rlabel metal1 10534 5202 10534 5202 0 net25
rlabel metal2 9246 4828 9246 4828 0 net26
rlabel metal1 6394 14586 6394 14586 0 net27
rlabel metal1 5007 15674 5007 15674 0 net28
rlabel metal1 6072 3162 6072 3162 0 net29
rlabel metal1 15456 9146 15456 9146 0 net3
rlabel metal1 3174 13838 3174 13838 0 net30
rlabel metal1 15502 3026 15502 3026 0 net31
rlabel metal1 13938 3434 13938 3434 0 net32
rlabel metal1 12006 6324 12006 6324 0 net33
rlabel metal2 15042 10948 15042 10948 0 net34
rlabel metal2 15318 7514 15318 7514 0 net35
rlabel metal1 14444 7446 14444 7446 0 net36
rlabel metal2 4370 15674 4370 15674 0 net37
rlabel metal1 4784 9486 4784 9486 0 net38
rlabel metal1 8740 8058 8740 8058 0 net39
rlabel metal1 12926 2414 12926 2414 0 net4
rlabel metal1 6808 7922 6808 7922 0 net40
rlabel metal1 8556 12750 8556 12750 0 net41
rlabel metal1 9154 12920 9154 12920 0 net42
rlabel metal1 12604 10234 12604 10234 0 net43
rlabel metal1 8694 11118 8694 11118 0 net44
rlabel metal2 6762 11866 6762 11866 0 net45
rlabel metal1 9522 8500 9522 8500 0 net46
rlabel metal1 9890 8568 9890 8568 0 net47
rlabel metal1 13984 12206 13984 12206 0 net48
rlabel metal1 10488 15470 10488 15470 0 net49
rlabel metal2 9890 2587 9890 2587 0 net5
rlabel metal1 6670 12818 6670 12818 0 net50
rlabel metal1 8280 6766 8280 6766 0 net51
rlabel metal1 10810 3060 10810 3060 0 net52
rlabel metal1 3220 5338 3220 5338 0 net53
rlabel metal1 12926 3162 12926 3162 0 net54
rlabel metal2 4646 9248 4646 9248 0 net55
rlabel metal1 7682 16626 7682 16626 0 net56
rlabel metal1 7918 15674 7918 15674 0 net57
rlabel metal2 12466 10778 12466 10778 0 net58
rlabel metal1 15226 9996 15226 9996 0 net59
rlabel metal2 3174 14348 3174 14348 0 net6
rlabel metal1 4646 6086 4646 6086 0 net60
rlabel metal1 15410 3638 15410 3638 0 net61
rlabel metal1 3726 3026 3726 3026 0 net62
rlabel metal1 3634 10098 3634 10098 0 net63
rlabel metal1 5106 6834 5106 6834 0 net64
rlabel metal1 3588 13294 3588 13294 0 net65
rlabel metal1 6394 14450 6394 14450 0 net66
rlabel metal2 2714 11441 2714 11441 0 net7
rlabel metal2 12742 11730 12742 11730 0 net8
rlabel metal1 12873 15470 12873 15470 0 net9
rlabel metal1 3726 4794 3726 4794 0 row\[0\].col\[0\].pe_inst.a_out_valid
rlabel metal1 6072 4250 6072 4250 0 row\[0\].col\[0\].pe_inst.b_out_valid
rlabel metal1 4002 3570 4002 3570 0 row\[0\].col\[0\].pe_inst.have_a
rlabel metal1 3772 4250 3772 4250 0 row\[0\].col\[0\].pe_inst.have_b
rlabel metal2 4554 8772 4554 8772 0 row\[0\].col\[1\].pe_inst.a_out_valid
rlabel metal2 8142 7718 8142 7718 0 row\[0\].col\[1\].pe_inst.b_out_valid
rlabel metal1 4232 6222 4232 6222 0 row\[0\].col\[1\].pe_inst.have_a
rlabel metal1 4186 6698 4186 6698 0 row\[0\].col\[1\].pe_inst.have_b
rlabel metal1 3818 12274 3818 12274 0 row\[0\].col\[2\].pe_inst.a_out_valid
rlabel metal2 6210 12036 6210 12036 0 row\[0\].col\[2\].pe_inst.b_out_valid
rlabel metal1 4232 8942 4232 8942 0 row\[0\].col\[2\].pe_inst.have_a
rlabel metal1 4462 10540 4462 10540 0 row\[0\].col\[2\].pe_inst.have_b
rlabel metal1 3726 15470 3726 15470 0 row\[0\].col\[3\].pe_inst.b_out_valid
rlabel metal1 3312 13158 3312 13158 0 row\[0\].col\[3\].pe_inst.have_a
rlabel metal2 4370 13056 4370 13056 0 row\[0\].col\[3\].pe_inst.have_b
rlabel metal1 8418 4114 8418 4114 0 row\[1\].col\[0\].pe_inst.a_out_valid
rlabel metal2 10718 4964 10718 4964 0 row\[1\].col\[0\].pe_inst.b_out_valid
rlabel metal1 7176 5202 7176 5202 0 row\[1\].col\[0\].pe_inst.have_a
rlabel via1 6486 5678 6486 5678 0 row\[1\].col\[0\].pe_inst.have_b
rlabel metal1 9108 10778 9108 10778 0 row\[1\].col\[1\].pe_inst.a_out_valid
rlabel metal1 11132 8058 11132 8058 0 row\[1\].col\[1\].pe_inst.b_out_valid
rlabel metal1 8418 8976 8418 8976 0 row\[1\].col\[1\].pe_inst.have_a
rlabel metal2 6762 6834 6762 6834 0 row\[1\].col\[1\].pe_inst.have_b
rlabel metal1 7038 14484 7038 14484 0 row\[1\].col\[2\].pe_inst.a_out_valid
rlabel metal1 9246 13362 9246 13362 0 row\[1\].col\[2\].pe_inst.b_out_valid
rlabel metal2 8234 11968 8234 11968 0 row\[1\].col\[2\].pe_inst.have_a
rlabel metal2 5474 12619 5474 12619 0 row\[1\].col\[2\].pe_inst.have_b
rlabel metal1 8372 15130 8372 15130 0 row\[1\].col\[3\].pe_inst.b_out_valid
rlabel metal2 5566 14144 5566 14144 0 row\[1\].col\[3\].pe_inst.have_a
rlabel metal1 5198 16218 5198 16218 0 row\[1\].col\[3\].pe_inst.have_b
rlabel metal1 11730 6222 11730 6222 0 row\[2\].col\[0\].pe_inst.a_out_valid
rlabel metal1 14536 4250 14536 4250 0 row\[2\].col\[0\].pe_inst.b_out_valid
rlabel metal1 11868 3502 11868 3502 0 row\[2\].col\[0\].pe_inst.have_a
rlabel metal1 11362 4250 11362 4250 0 row\[2\].col\[0\].pe_inst.have_b
rlabel metal1 11730 10098 11730 10098 0 row\[2\].col\[1\].pe_inst.a_out_valid
rlabel metal2 14490 8806 14490 8806 0 row\[2\].col\[1\].pe_inst.b_out_valid
rlabel metal1 11868 6970 11868 6970 0 row\[2\].col\[1\].pe_inst.have_a
rlabel metal1 11178 8262 11178 8262 0 row\[2\].col\[1\].pe_inst.have_b
rlabel metal1 10672 13906 10672 13906 0 row\[2\].col\[2\].pe_inst.a_out_valid
rlabel metal1 12972 12342 12972 12342 0 row\[2\].col\[2\].pe_inst.b_out_valid
rlabel metal1 11638 11186 11638 11186 0 row\[2\].col\[2\].pe_inst.have_a
rlabel metal1 10396 12614 10396 12614 0 row\[2\].col\[2\].pe_inst.have_b
rlabel metal1 13110 15674 13110 15674 0 row\[2\].col\[3\].pe_inst.b_out_valid
rlabel metal1 11638 14348 11638 14348 0 row\[2\].col\[3\].pe_inst.have_a
rlabel metal1 10580 16218 10580 16218 0 row\[2\].col\[3\].pe_inst.have_b
rlabel metal1 15364 5338 15364 5338 0 row\[3\].col\[0\].pe_inst.a_out_valid
rlabel metal1 14996 2822 14996 2822 0 row\[3\].col\[0\].pe_inst.have_a
rlabel metal2 13938 3859 13938 3859 0 row\[3\].col\[0\].pe_inst.have_b
rlabel metal2 15134 10132 15134 10132 0 row\[3\].col\[1\].pe_inst.a_out_valid
rlabel metal1 14536 7990 14536 7990 0 row\[3\].col\[1\].pe_inst.have_a
rlabel metal1 13570 9112 13570 9112 0 row\[3\].col\[1\].pe_inst.have_b
rlabel metal1 15318 13838 15318 13838 0 row\[3\].col\[2\].pe_inst.a_out_valid
rlabel metal1 13662 11152 13662 11152 0 row\[3\].col\[2\].pe_inst.have_a
rlabel metal1 14260 12818 14260 12818 0 row\[3\].col\[2\].pe_inst.have_b
rlabel metal1 13570 14416 13570 14416 0 row\[3\].col\[3\].pe_inst.have_a
rlabel metal1 13248 14382 13248 14382 0 row\[3\].col\[3\].pe_inst.have_b
rlabel metal1 15824 8874 15824 8874 0 rst_n
<< properties >>
string FIXED_BBOX 0 0 17202 19346
<< end >>
